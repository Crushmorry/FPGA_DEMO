

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EhEutCv9KlTIFuVGm+vsqpOvTBpo12RE/p/1ZLq6OJuSzv0CX5JVucDsO8HJjZ5n1scocvuhrD3v
43PtdSZrXQ==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SH3/bIYS4p8YYaXMrIdzNE7Fr9HSHFi38/v+Yunc6fPs74Z9txPvtuKwPYj9F2RGcvYIFjRbKWfm
WT4bs++O44siibKqmQQNWxm1Sk0CvlqM9wW/4Q7VLemjxEL8jKqO7RlliaPx9dyj2tLZtNyZWYcz
Z9OP8+MdsYnfqU+YgL0=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0kdhclGIp+Fl8WySR1hebHNshSQ+yNZbxYvclUjJ7+0WHPQxZqeEZ/tcgWpjczzWd+4OAPo/9HCc
X6d6SdcV2d7qcgIGc2OOjEO/aKNKTadPONuLcB1qfiVG3He8KkDmIZUZ8fIyXc8Zttpex1HVD1fx
ymY5qSLQnld0SJdx6E3/oja6P9m/26/cpp1HGF2zgfluXk+sl3nfTNP/QM/HqEObWL/MJn2K0st3
5IQMCxinQZ6vXtFusIoNXHP+HxHZgC+MdrqwCix/sg4nLZ3iOnInSo+fSdhCk6ndHI/VGlTAq/tw
6OjTmtAzAHPPmgHUc7TFkd3dyEgtKMKb/YBW5g==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
pzydioiu17Wl1dUKNc9MCpMyYzLve3DG1DipSowwELFIdgdHY7mGykyxxRJx0VQ0P8cbE7Y3pNl+
0/uqforAU3pGnqtK1d/7fIKO/Lmex3YXHfibZVf486TO+g0jcNAFsm4yJBEAemUfgZlMtSBNv38j
vHNdaaBsjHt2r+Sry8lg8xCHERRX0H9A+/ezVrUoTy8ETLJ2wyoSZxQTPadf/f1E06r9lrTmT3Gv
HpVQRozlNiMc8ublXnABGN3UWzVUL7KhVSQbD+dfrAv5SXZMqkT4HYoyqlHiLJd8C2p59wnJqbNx
j1MZIsLW4ZpphYsus6NnuMMAOuCcrU5ne+xU4g==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
YQdKtXxGjJdELkZmx5IzWvetY/pijiGXvMWVhkjcjdGj9WfZ6tCphc1Myyaz7laC7ZpjtZGBmkB9
d4fK5e0+l4BKhgCRtzjfQjPN+6cYo8Vq2ld4TC5NNew+vCF54JmtdG/GQgANBVhzmp/o/F2Rn1Qd
X8LUj5XON/ybg7NF1Kc=


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cQ93Y5m9f5pYlChIpfvgQ1eW9gwohiXhKyaoXBJiUkkhdAShCtwI16jBxg0l9VHAL0tc+ifqY3jV
jtjL2vF4W39a6igkp5LeDA1gvqb5yxgSM7hmHjstWeL0pi8VOS6J98X525Zm+q9wCXtBlpDfsG+Y
9YzK+uAzUIDI/OCkpMZCc4Opk+SmcGY14H91ZP4iE2qauNja9pZYkoT1dljIDmdbp0HoJM7RTglS
YrMH1z0fz7wdnTrv+F1BqX+BnMH9mYonM5mXoCrVvBBQUoieYwVfLuSmlE4dI+zlPep1IJgpU6o6
9XrDEraA5w3ob+eNKT5Q6p3ajAuahyI7Fh6Vnw==


`protect key_keyowner = "Real Intent", key_keyname= "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
FEWh/VHO7WtKkVfKnspXfU+JEGIHgTbsQNZyPC/uBHUTkmRG5QXkhc0DaiyEm1GWAXvcNVxqYLFQ
sys4RChAQLUIL4xtXJEC6WQQEx3bNXmlN8zQVWTzkobJiHRXmLakzTBlG3WKcJf86LoKp5l49z2X
OMUn04nNN6W58TXSLyznPAZ4AEuDQXoLxbeMwFV8tca5vsFii2hqRzTXgbsywFy2y4B9E2+lfBt9
SYnvM/GcKV4EmduTysSUzN3rXYmyhYZY22VPZK+p16UW0r1rgxbMvg0Dv2z1tvYXCxCTy/ncEz5e
zp1F6/oLY9LrdL4RI9U8m2vlag5NiyznYnKscA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2019_11", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Z00vSUT4j8kxSO7Y8k0hDTnYto0zcVHNByVUFk6GlcOTtYIenU+8sIqapy5eML2G3ujMHQmlf/zK
OCQ6nUyQYbt5ukdvBjhJ2mX+EjC5HyuHBeSf1pfKN/TWYwPxFGX+BmiJsxDZ/a7RFE+SvCsLvraj
coCC+BjPJvEp7fdVFKkkkklqzimfDiOVIW+ecacV7yplEnB5nMCkF4W4wAu/Vika0KOnzHhDX7iG
ZUkPpbkYmlMXEs4wcBeYXRrK02T89OLz3SWlbDhodT918Li/KEiCM0VXP0PP44wvzAe13q7jvpwm
TBj3KdaRuQ2bezRjz34mkbCG8hwO+CS49mtR9A==


`protect key_keyowner = "Metrics Technologies Inc.", key_keyname= "DSim", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
YAi0AO7tvimsyndmDqt0Pd5dhk/ZmzfDr60rh6gIOwktCdqnn5BpXmteSFkoYk6zBgRIIj6mw+qB
06UvLf1W1jXFDQNnRViq/66aBpEC2Cir5HpMU8ruiS2rXY7GbdHTFrBtTz0iCF8m+StXYf6WdtkL
/l8U7W9c9UPdAovUv7CFb8N14eAA3mksobhxpdYNo3P5oRQ2/pksJxisCQSTQ0PnPMDQ9OZk+xZk
L+jnGUikOQU3GcyPC16dV0LZt30Z/pGStYk0VVL9MTg+lJKo0ng+iRw0un9CikDflJdR02bdcHKb
Lkq2OTyHgPfJO7OPMbSswzHdNwdiB0qy6y1kog==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 334096)
`protect data_block
D68taA1tqE3poShajgismzsmtd/X7SC0b2dglmoix0rbyJnJj7m2dEdErqb9pAQKan/5TGQNsdxl
NM5jEXst5NVJHYloWRe2UqTLOA+k0HURMzT1eDHhUOQOqdz33rhW30FKWMpoS7Xy6V6jVUcdCC5y
42dn+Vju5VMiCFRaEsI2M4gWBthpWzI4ASUvUkuj5Ivja36oJRebAE7imvmhX8TQ4U/wDl4BwMVn
CxYkzA0Lcg3GYsUPcsHceIxciUnasFXdCR6g7sGmU6KQ2/05cTfbEcvVfgMmX7X1+zQ4qjFED4ip
le5iTyEMGz/NqWcbIPe2DYXhd8n5A6N8lCNgGtO322CenGJvckKrFu4rQmxLwZ+dj4mOGNCQCS+W
8qXBhgn7FsLIJpVeiyocyY0QchG4eJ3FnyeFs5x4sQfbbxckbhC13tFR2n6hSen6obhYBM/koiEh
JjVxJK0SE5FZ5uYCMHps9LLu5EFdc5fmzsMZ0Q11QZDCI+UfavnXmo1R6eGgvaMmMpB0ueZ3tP4t
e0lU2QQ17QuuIDab97KJiZ2bqVW9E6PQN/+1RYIwg0GtuA7ZQbf4NhDVY5LcaJ9WgE12QqyAD0ib
rvALpZI/thYXIZOsL41zYVPPI1dU7Y16uVIF/5fe1Keoh6D20iAjMI+phmlt+7NfMQK5kjJjW3TZ
ciXTpcRgqMHPHV7OmyOtHNwRB/oGJusE13eK0v1drtIOCfIlqUUqvjiddjs8zXC/eQXliAq0PXEe
JfxxmxTnLDg6flLXZRIodlN/an/wUqbFV7R9gRdq+KCg4+YrsOT0+tU3fwCuQW+52b8Ji8aOZuWm
7/DL37GPN2/qvf4uVKfmRsqIVLG7qxBb0GXhiQV+wvch5JveGva0B3c2FyLG6mGFS/8+/fo+5s1E
4EjzH2e6sBqxJQtHO0fOR1fNx/Qtqfa/8jwoqnniMz9jlPNkrKanOPPq9vlWTnBJ6UJDFEOuhrtF
mYAWnO9+un+CQW9ytdXrJM+xhKAVHqyenHXFsTrhHjkhcio5i5oq3Y9I/jFJo8vgRfR7jgegqwQC
2rLufDOEzvRgddFDo8IzkQETZknRjwOza1oVII8kOi47MBM3qjD32xAXRdHpjxOcaNI+ecVxsTVW
nwuvAo9UlA5sOGX7kNFqcUK+WAXyUOwBgwnQlbQrWBP5kfWRSeshU8vQpOcZ+Hv/0BTASQzfEvBW
dTfaLyrUiwKfs5YSnyk4crG4g7ahji73Z5heVJeJ1ZkJzaTDhcyizvfQFJITM5aqlq723mS0kwmA
gLHhz1iBwHNoyjDpfLnr0b7e9AD7cu/mojVE4IUZYaxNtDyLd/9EMihXiDwj2p6fmrZiX5+A1Nhj
kteVK/sC8WQtOxOmtoPd5C85JuYDOt/qh32PPkFad17HNp5+lpd3wvZ2CUf4Y4Twa9IUgCAUcyP6
qea7yjl06NKUQhFor/OZ2MCNWcCF1HFz+8REHgZnmAvEd0n8P8BHf9O28YCZFy/RkJqzJiN3ypW4
Wv5GjJIgKt184/KhtOSKqaGRf9zJPciSbx+LPc0okbroQAZjBw/ERgjTRk8Nn4VhExItd6pndvy6
1ADAONyhkRGFDPnSQWd21i7ZzNcGM7ItAWrK26/0NYzbOenP1P7DkQ8Eg92OE7ZfXNVYMNeKViSY
isIcYZFac2I0bwOj9eC1YpPtmqeuXRaKALv+am45jMAvk9cg+McEA7afd/PWmzTSnihqVdrmTXgj
PQcUt48HFs6dHJYa+GbkBvynnHnh5ckKEmAhNo2maZ9kvBVekdxCCHrOD7T1jXN/+U3nB9CigXH4
M92nFdN03aRlCfgAkfQrui117vNJH88XyN0b+qOUsbyQocqp/WJA2g8dIY6Ms0RvCOWrTj2aKyap
21AaZYdzXUoVx+Y/5eAXLZLgcC/EIPI7eDOT+u2oOYurcfO8lwEPhAjoiOkepklQaBwLG98ERcCG
sZshp9ADNOcjXFwMo6GoC2kMEConuKQ4bRTZzmKYQ6fz2FnEFsd/jKa8wdQj3iKIQQH0aOOon25x
CUuFRP3r89xTsOO0yy+zQAYACjFOxfhOGf3Nlr+kMaMDiiOrPKr6MnyAYcHNEgqzopebanwtrsa6
vM/25aWDwyIU6j4fmXCHoPXywfrW18hrx2Kne/Lqc3qQYZ/ArQwU5LkDuOC/bvLRsoukgIU8bhS4
DUDdw/TEiqh9dt/+bCYon1UCzDXId2eYPRXS7LLli3Xc1x8wJpSlFR9k/OXKyMWa2Pq7mJigGq27
ndxCCGLXEuCxQADh9gpTi9SzOvhQfh6ygn2Gv5SbdNh/LVvTbLUiUku52t6VDXTu02qeDW1EWb/E
KrfnKVu8wJo7SD9vpORsfmCBZercSz5wtb0eIXGOh718pQRAVX84DPj/wav/Rw9zvEfg4nIWeUpq
ADRaDO3tdaGz7RhApf19GRQC0cv0n6PkdnxnHCdk54Zv6yPD0mKV7FhjaSSjq9p/vRXz3cD6MbbF
hlwQ8+0srgo9gmChPplqhTFc2pbYXbPNhxzZXlaV7rYeF9cuRGSMjxWyz56VG4b7cZQeCumoPh8j
tM2Mios44jYfp8nYm/VjpGPU2vUQTCbVc4l7uY1M76h2UIx409xYWF4VjPT+eC71GXMDLGrXMBhG
vpT1XVbeQa+6rxcA0B5hYl6xVoHQdwoNR5Dhd1keF2ENK99OxPMxkFbM7xr2t0Iiv8XvsMasqFUG
rvnM0/pHChdvLyjziE2dUejrpaPxKr0HWVkpt+57YCzhCXlAKwbUnpv0xjtpuFAiq2DGeVtGSgEN
yPavyILInojTuvYSim4OmJTpokzNgC4lm04AwnMpVICFEJeGPdjYHXF48oaJNCA6xTLniRdWyaUi
s+OIsLLxlYYxDqnldyLVJosH3xCna8jJ2CckgLylWDX8/Q2Jv1GCz+0I99oC7lNVJeXWE/BEFbJq
Ux3XMuqdmR5D3v7fc6LttHp6HJooy0feOhBp98Ju3tb2G4Scev/WCstJJ2AncjkZlC9wYi013AsF
n61zY/lrouJQVlI5UIwk8z+49hBYkY+LlSpSCrd2EYUW6K3Fm0+sROaVRCQAMlZDGpzYwdpVs3K3
BNTaaOYxAjgQJAHoB/hGSWjwOYg88Cs84O/mEk79NWWX5xm2tlWW0Qc1MwFrkLaJwmB3MIquou2o
/EGgh1KpUvUJxJ6zMA2BonB9RHgZiF9GzCibeTpdjzo9Ke4fFw1Y4hVFVFgQXSV+bdZb4/NG7eIO
bdy3cNk0T5YobqEqBgGi9j5/ZtNuEFXoviLTe/xABI9SGa2/NQPST+Pb0VXORMpRtiGAWIJiJz4o
+2egDncJk4glTWmZtRcGEQxtd5FFcCPIRCRerV7KbYfZQevZiAImI0ctoEwCZZsLj52fMk21S2p4
UIBfz6zA6zWtUaubuSMccXq0lY6lm/qyPznTbTGFCYln9AOsfi0IrjWlaS8Lz/XHVC53mGJEErI+
3Gia2BRobwmE79GKlL2svmkTHtJIF/zolnsEkj8CmGk3/T+Wsd1TCM+Uon6vlwc4qF/aa1h6F+38
lKlEIdxRb7SPIiqfJNPWDyq7mYWWaBWLw57xBR8dhUJmkY7OMGqOYG31bAfmUaKdlCNQxv29Exv0
ZkDGDa1KDOaQY1JLVZYRmryKzLgQfLlcR8+gMGxB4KHuUnyPmACvpywheVL/4gS+sKqinkHaYN2F
2+ymAnBMQ4Ug3sbWLpAvs+szNk/dJcc2JnoymmVVBAoq3ZJysm5vrG2yPBjBgs1u6HPZfnr4TKgi
vcWakFSkK0VVKxLIs3LZDicBxeAg5jvDe/ACp7GbNnf7BfdIHSzhXxJXF2KUNCalffQ5dTObnjG+
qd53VvMX8W3zlCy6xE40OG/a6GhiJEimaDkXr6KBkBxRGXJotWu8e9ct1x+J3q3/j3pXRsSoYDh3
MQlnO8KOATbvp1e18LPBh5GO4oGiRr202Gr28knz6bwB3uHwAAsqvGWB5JGALVGcevNPnEBz++kZ
6fYdquG2Qukeg1cMJ+m7aXZpWRkDbz0LRyrIbI8ZeCkX/k/juB7Vu47IJv1cl3FjTLC1HUeb7TIh
tgcb75CNcALAV+DInPfYNAHrMxJ+ikT6MCdWugU4ZHY/3wUN3YMuVYANTT7qENhMIeRRx019QARb
RwavBfGAhcmj4YCgjeeFswChbyXR4SultcwYx6Y3HnJsK/nCA5aZG/eNU2JqDwbjC7s6bt2keY6u
7PiZELRwxA4r4nwzLTgvnH7ZBTYmSZ9Xe1pEtw2aIdO2OFfG2NdAq16Di33tlJh59VgY9phDAWdw
3WXxzASKe0s0kFRxU+Zbbm60yO6IGNbbYGGhqjpiKUUMQcQBm4EViBobd/+lTh/+Kn5munlIM2RM
WSwQoM/l9A81Rn0YGRqJSwTAmCooIoRU8LnCmECGyspHcAYh6HtYbpbaeU0oML079Rbi+9uVbbt1
lB7jm8531bCD3bYwrBarnuTOJTefdrQQgABtAMCZ7dA8K31mlfiQ5riLHLehtUVYBU22/7QhCjp7
8oQ/vb2Qu2+jPykPzBfjg0/P7sPvXcXAgn0zA4O7vpVhDjgW1WB5vWnIouPPL8cnWbD1DUK1A/WU
Y5lztMgELaXK8JFAyjeSgFnSS/VKrVrYj0ZoxA9W724aFtpzRmklbN2XdRWr9gxw2WklZTa0cMnB
qzeTnhWuq9WaOucWEJcyR1kin8WqlbzOpoX11fzvTKX6LfctxOMevd5FUnZwv1JyyW/5/AhYgBji
/8H/UwICLJZEUilzMX5C62NbHz1yRsTWzyOr8x8mBScIJqaFLWzXDlCtKINA4w3InjRfmBioWeSH
ZwAa9dyOPqR6oSxCPWIkcP0pUqK02KotBeGZQm1hytQd8QuxQYiC8wQb+Y8+4T+8IqEOzIGqfW62
iTf6xT9aNQU3rodTEEC/L85tpiC4VMrH44robg4ZZ4xh//2bnYYVTyZ1OiRozPWF+PzHWICwv/4l
DFIOqZYTwERzBVlAJhXgTQjwZHykLzqfQhFOF+HYEIFPPAjPTnA/UZTHX1Ltefn0OzmRXgYj73CW
90UV9Z6Wv/p7QbJFMzu1tJ1BKCFpq0MIOYqhF78RLeCfPHjn3/TOW9LMvPgDOVqz2KWwOXLO8PRd
9jjNx5IRM1uIIqNfpFCUhC1xv+3foUpDilVOSkuOMGjRP0tcKXuAUfu2Jur6L5u7aymdrzB90kXk
ItFuykOHAHK2BzZnqSyp2DWV66GdUWlxCWKSEDfiMigRDCpA+jZQcy4rfdcEi/vVZDgWEh/yEF3e
2QRNaTMl8WIhW7LHR/7SfTX5c/R387BSlmT1naZzpgCqjzbJpid9M4k51EGKsKRH0zHCbefvsKUR
kQdXT3SaQL9YZ7i2kuiV9O0aBfMo8ivWCHaF9oeF6JeT/eDgUCoKt8vgo4F3mg/00Xx2+hc/FVAY
bM0gl2szpoxrYpAm2CD476BGVoonN16SQUoGQHtFf0aTd2FTWU9Cjyn7AvxzFVgJzwrm/0b2OXUM
caWiAoyWgeF5JZJU7zhu8Co4F+UFKoS08EDVoh4GYmozWoBIKXouHvw/YyTYfpex17xnQ1QXPmiC
Q+k2Po21K6uy4LGPIIAjthioeTUYx/MHwWAq0fDoDB2MdTayxc8oV9lE9+0EuYN+84KDTZuZyAm+
Mrhto9ArgwnInpFhWKIfPRrdTDpR9+kO/eex3vcJE8WaxN/+/P8r3NwljP25pHxFKlS9GaGCNzhP
niBbG3ar7a2VHxXuCh+warVvwMF35fX1FYMoFNEbHhnmaxvKjwPtTz8ZGMZ4Cf27LKr8+wCzRs61
4VEdVh/VTJulFsvIu0nM1YKIlNuKQcY/qbNe7YmgkskPcUCAG33vanAtHjbF/Xcmd8kRdJuU1B0z
mipK9TiVdH5XDzf2uNrwrO7+Kfd44T67X2BdistpGBJCzkiizTMp8mcDlL4LbmnO3MKFFEDImBfi
lm51hPuEuIF3EKbnb1xLTE48p8s/qST3TOOKRDq/Dbo6iuOkgRe5q1cVS6XLVPUMJlZCTu66YVdL
moPTWYhIjlPfchJ2Eek6MzgdZM3ZnQMiusx7PTaSUtaWZOIHmUgfaR7hClowdCa8A8+KAhjLyMIj
7377Z+Q4rPKeRuaExKdZ0fs7urTARMjxQJ5JdT//TLxMw7NyhhSVFxF+0vGtFJ4asInZdtjDvM3S
ZGNqJPVBkTrlxvITfa4pT8jRrwO+V7h+LqxT5U+w0np9T1T2onFg9fwAok0k6Fgayz88NJ6kA7hr
t4qdSa/WLomuOGOcve96mm2t4e5h1d7UIxoa7+d8mG9hoqcoYKi4PsHGIM2OoZtrnGPCVMP9YmBn
JKhQGQrZN9W/lHSyNMd8lPjbepog0aLnBwbrZX+u6XGYlBWp7Gx432FFGmvHSGaazIvswslDyFxW
DjR8SO7KWHYdBT38SpeGVn/zSz2sLF1h8bhZCn+hxVso75VRak4iokyPcMaMjoDj4WvryqgSvOSK
o+A41MHIyEKAV1t86j04SrJDY2RD5TY3QVFzxCk892NjUaOWxV0Z+CTlo2WI7lJ4o2+7xwR+yR57
rN9iBqUPTfHpVUnGsUqS3JNwrFQP8t2NtXtBi/8APYfheHpf4NpLTWXq8lmMhasLWRJiVhpKeJP8
Hll4eHKXxXYhGR6QO9+PhsgeAGtL1uQN/UhM/TqlrT+ewaV5gZYmghgsIr7oa7YBATDAie3UBwKt
4swuslfGJ+PNXf+PfgL65w16vVb3KVoBsVwyX9GQsP1xo0OAmEJPFV3naQrt1uE8KnfEtMMkaG0u
xcZCWLIqHPyAapfsD76pSPahNB59MJhQwWtqkpkoBN41LQM2kUNdTKKN6CHVP/OH1CXht+H0Xlon
MtEVC4MVUn8Sfmilk+BSSiZlVqtkRO5UTa+wxg8R3C+t2A1pixUiWG7FihQwCYDfL+wD75h8hbt6
QQ8QHQ7CNEM1Z6pjgYd1BmMHg/RNdgv5o0zo7P64cqBD/YWv6g4amNwnPYvyQCw+sfKPxVyVc9FL
kHhH0/leyEJUyAPpOr6r1/iMOPzyAOalcarL6+HOhdNEHQCO9mCR7KO9QQrxWmvxHLGNRTdLuIqF
93TI14CCE1giTFCxRzqzsHeOH76zs6dWIoeDY8aPl1VuobqmKQZ7vymDgNY+FrBaeOkQQA8ETSD5
Y5Ar5OKiHMFNX4J0kBn1w/KmQ5Kl2357CBohy/TYvHBislsE3seFLJPzWZfkCRVu0X/Eyu3KMLAS
X1Am3oP8SDDcZfx4OEIWnVulChObeGnepH+WqAylrovZL9rf8Z5iNI4bx/mWXc4U5iG4inz1Eh3i
9dZz/upYwhgbcEPgs6DYc7JoN4KH1n3ra9PgQH8Upez82vew6WtFkySh/1rILdZHjDFyuJFWBTTz
5fIiegS+nuqE0NDx71iHhHLF2WNAyDqV15C71oxNPjGP1kyIMyvJYog7pHqZNeXQBOEExDNq5qEv
05tLY8iKF+CgQXAfOClFI+4DEG+d7ga+jYvKT8Dl2D17TqkVvG7lYSDpwL9zulILZtXiLN6BW2jy
mblT0jHiBcR5Jav0BveAHmzo4VQiZPF5yneO3I7o1xaFjqMWmzSFiyZKI12lyuBgvd6Ielv5cp80
u2c1aPFE3JIed1FtVP4dk2ZFjOonRFSHGyv3mQH0NmK5AazLYVKfHeRLwiK2OBj8azfr9T1anm0v
gqkYPEBa147FTa6WyH7Mx1vaiMyYnzrpECsYCxb4hmgwRgsH3NUae6eN3GJuwJQN8GCjNt6IhjEb
qeZIh6L7BEcNgneDD9cRCvv4a3yeM5iq+kSd26hNRB/mxrjXv2w34MxlzMeB4zOwjkaAlkCHLP3R
Hp/Wn9JiIL8MQIDO8H6FpqR9WP0TNtrZ/FDUhmfKjPkBPftEljqKe2KExUVGGGsgUjejc+vr2jvw
67GYiGzLgJpYjrYkazfJwzy+htF8lsIM/XV2LnrSqxpOV6zo/VWMUnyraledXucEAY/T4Z2u3n5f
xADG2roIayMcmFX/TWOgp80NL5iDyiSHaO9XMuDrnOWOuaCPbpLoMn25Zfwa4cy/Ze0Unp4wvFVh
fQvfY3W8wnqwY2y9X/tDSVfoR12MyU084yYDfjthZa8NOaHn2+z34a/1cjD7urLra8Z9bDC5gtfs
hO1I5FcGUuZ65xRXYBXwPtedQJEdZhPKiH0DyRhRksxJUYNP5gpTt40/EOrA00es+LnfVnauNoxI
uFPmvR+b6b+1vI+REDkbzm7eZqpaQiTwUKhGw/8T9q8OKkbgjvMZoelK3VUx3z13ruHVzyeRurEw
GQgajhfsuWdjBGklMKQwvLhC4YKW1qnqr/qT/dR7QqTCUKD0yN4c9KSdot6URsT9o3qkcs24Y16o
Tks60J+SLMxdWRTJ3E17XXlp+Y3TJVKNnvCstZ7NvwoNl9KUJE7e7sh5D+AyVaW7UTefG/q8B3Ov
fvxUoORSVvjtMOENLKWWjjhLgyqoj+iNI/yJiMtOl2oLcO114SBpYQo3oZ+wT7+EIdldTYv4OuTj
IfbJbd7ABFHELOHApu9Xwda6hdik63XuCaMM8bpnZi00S12XkDyAm9SOCdSVmFhY0D7s9Twu9qyP
zI+4uk8oolCNrF4CXJCZOZ7hocUN06EpospL60BE/Tq4hcqrijIcmxCd+eARdBO9Md2cku4wztxm
1ZN960REoQDUnonradxK1pllGF+CBY6p+VUXQH8mlljQupSfBdkiNVGUMl4NGHZIHZd6ihGi7a+E
JOwQQ9NkEwSoICIzOiQY3STtQCns2ZiA4/vjIJQBBc+jEyawh1grRjHgSHQFPugzS+ZL58LGwGFX
yWYSNvmTwUPIJRYpfzuY3ViWy0o87VeSMkH+K+MCJu8DbC6pVv9Y17i6LZ71cWgBh3sZAawGerKw
5CM0DFswJTKrSfogj3PBlclv4XOwC7jsT3rXP2oi5Krx4So/awF1z3irNnMCG8flC15zRU9j1bqk
HvTtKHg3GaK4mSNwp+i8boiBG93dOWMg+u96huUk+fajqRYYlU4P8lxc2+pWRgz4uIiVjqY6/Ad8
n2znmUuw4B4SDBKbUqFXNoXetfHC6c3tCSamD/gro3au8h4BPviS+9d5ItLYZxhIclQniuG2E/MR
DZ5hb3pFUV/Xntm8e+H8RwhxmIZ1hpPuDIVluTDzwyLjRvOZiD2TH3nMNzz8ETYH4m6tFhYe3NK6
x8/krNkRJRxYQvf4UP7q59hqrqQ3m0DHqXfUIlrWnq4XDLPXUSVlvGCiGpELntMpbBlxSHgAwB05
o19/qwoMRNJ+asXmQibuwwW5SnZxqSEVMnW3Ov/acaRc+57/3l3ut2nGlApWbXQJlIn/+t/d/TYU
XLgxM7nLNakTDD4m9CiZXOxM8vdJ/CzHKoIdp6nyWDE0v7CIpJN+hAResu6skzm5Fpa+TgsKKdkK
qXGXsqHkPTGj90mTS0lw5Gp/o65CDyaKjp0xFXgX9DhkC7Biiu4t+AnW6d/iTbKXRMyOqZE4AabR
MSBsD6Nrs50/ZCYPnmCLuHvi5HGFeEnNX1T7kqySUAT2385etNXuH59pJVU8TyZ3e0L5FSj98Pw2
P9JAX4ZggDOW7ti4DTt6OBWY8D1s4PMueBIQFJH2BzWqxfbGWHz5OHAcn/ly+cCDOPnsGuNqK954
HxYcIzPzoBc/DApFYry3bMcMoIxbjKzYFgoeWesQOOZgKh3/ByRey2ytlO3NYwdkRKKvL/Eyamtr
jCFD9fu60mrPNhwXc/wZjz7ptkiwnIYyQSUmdM1Smx0g9PkD2CICn+BUb8MOdRLGJ3pN+cy5Yrr3
Nkp2LdUlfcXcQboKO1Sbz0ZRdNH8t/ph3dWWP7I3UDrm2sdAn/ro0blqKR8EwB4f4QO5HqFCzTu4
AY8iaqGlY1Nw1lu9zItHiU7xWEH4/4rqCCXLPhfmGXCltdYTJTtD13bODjGNqXd4/vkT1wix6F2U
ByrrFCJEnDwccZWHkuFwyEqxjuKI1rarz5B2l6234sJCHz54aiV2uxGiITN77+90oPVANMJ7Z2SH
0ZRN5qNNabXD61BTMwCSoTyzElp2sRmGfpTdoTdR50AFRe3lTcm2PrbhniZkVW60Drtx1gDmvsR0
hXmcy9KMQIIb57xOVzh6gUNCsCGFt1VFdNFtaa/vYSUHmLZAan8KlmfKtLT07rNAJyHrKzRZE2bx
9xZYi3w7Xa+UT+RFbl2v/tY67b1KgTPjTi7C2mBD9qVRAosmgir6htuBKN3WxT1zvv1SSBSHGHo7
+xttHJAZ71LZ3uEUgn8Ngqgf4MjLoMq/cv8Ell/bm/pZistR6x1IvcIW/9zV+5AlVAs74cHRQYGQ
b6anjMQzibUhpcA+HkQIAGjII1vgT3HQkp48h8hc/ST3BNrqUfSvykAil4M/Lfl9jf44N0OWCwgA
dc3l1AcFu7fqOmoaKJqZ8UK/HdY7WgiQGbte5L9dkW7uRNI4JI1HpJN4vOwO6kx6FqJKRPwtGGmQ
TTek9YwSITuNlbGpsRl9GVEa3Et8148OLANn/Qu7G0XmVf/gEOkcjC80neWrxyZFDyc6HQR8aWh1
9rb85gkor7skDW3TOrCPPUK5vZuEEwLlksLOuctOMZLy2/mHsiIt6r+vjubJ7EILrtcUrr/A/qgQ
IXk3eUwjs5NKSMOsCueX1zEfxBBZi5+KYxWfS87fTsgy8UnnED05MQm7tl3vpZxVpp11rccVP4RM
Ib5GIJbLOyPiCkHaLy9/XSHfMzo0hyM7o/iHN1z0G2ssHht1Enn6H0qzmqlh4DCTsapv7I18zIdK
16vXylt7K54Lp32Qm/aiB7UBarbSZSBEve0bq6AihqjRZYHoON5rpiJ/Mgq1TgDdt4zAXo3Xe/ZK
g6ORADuzMNQoO9NGdY5MAtyudyTKq48wnnoI5K1PJpF/8Pfvi0dStEAff4bmIMHU08UCYFYU0/rz
cWqAsIpSw4K/JnLHGi4dcnWuEcS3jZZfiWxSrvpg5iJ9tn9kYCXWv99idBtC10bF5sfQfHdGeTkt
zBRPqaGJgYK0bKCGmZngq/X9EOK62P2ndTcsZ6y5+iCd/ujGloLKHACiQ6Up1I9g1Qwrcg5jg5Wd
qG+1spJgxBgaAw9bK/iujF9rpMn9XBES4yCI39f1RVebzq4T6PppdptU+ERFyNRBV2npbb5CqgBz
IvhMWU6tUvnoiWFoZ4zz3ykclqdzDS/jW0bnB+qXn2Oou57n/HQwRw/d/rqRTnTKNcC6GrRSt40d
ejd14ky4Ke9Rr206IGSYidDYMYdaPunyvutVXOdPqYrmOquj98Ls8uSKRCUhJFtG4GE1Wn1z0EmI
krSshZ7XfIxOR6nV/BQWpBcdGbFpeLK5vQ2/YEIpv99WPi1k+3y2yusi/w3vD/s9qfzYMUt+3Spl
m/Hh1I96sEc/bjaqJfMY1/ahS6kZg/FUMReNIQjY0jHPI2TjBu6aMsBARwqxRoQcabDgdUBemFr0
8PTURapxktc7JRo9modcugXopaw4/T1xpxVZ/ufklxmJMAbfL5NG8ipi71gbxwWIKLJbuog8SMPj
RKW/yw3nMWU+9RP+f9bAYMKqlP8PtLUq2P55Hvj5e+ev1RI3AVuDgary0YwPPzoDKx0xK4OCeWNf
6+quGvW0vPo+7w4qR1H7qzVAlSLDlzH187On3o4WkcEN3hUAOBdOi+W1xecYfVLj89vW3Nr+6t+B
hfsKXXtMnI7CZGUTv8EsgFwWyOtAn1IshOp05USpkU5ObSxlAHG0E25y9zlmBm+bPRlCSFq8Vwk/
P198GcczyJWL0JGu9JCSuvYhCscqna57cJMQ6PGeyWiJHfbgEEQS6+3AXHWIVPvFJgjTpgCEZind
Z2gqkuJnIymF+Jvi1wHUdyh7N5UkVt73r2WKw8Gj5cscAbSG65nfhGnkk54fTNMxeCDwBVxoYUwM
zDPqe/hRtpHS3LP9hT7U2R8ZtIdA52IaW5oOTrTlXXGqfz6M2HCFtihMHSCfjx6lyUCjGb9qSCjv
am2vrpoaQwvtVSLVemL727CLUbkxQ7yR9lrazXiBL82foNZeG9qAjH9Z2HTR+JKsYIHgKiorW0Ri
T9f5196449XLE7ftMNKZgHCqmr7yDWs9l0G7qATCaDJYL3Ub3cHPLkTHplCm8AtD33BHBFpduKDp
wMbGR+2R5tBO7em5YInZ10bFFHZhykjhlgxAHv1D7pFmczWlMhDpTyd7Go4KvCeUBh7zw9OWOyCR
AS3FW4PBhnjqLauT3D7pK+6QcsWbK3+IHdTo31CKxMf8YypjWFYSFcUDhVcNZlYcuSjrwN8+fdla
5Gen4Lci8IFTJz7RCBrUcBNUuQbkNd3OsJYxRMp5NaE1C6+HIiek8OJoFw7fB1FCTeJI3uptawj0
ofo8YDS/QxXf8YFIgQbFQCDPI91rUN0l1/ETDe5sVFtdoB0xFQ/Z5Qt/8rwcR5mmng6w2uGMa7mN
GIcL4SYkzP9IQ8GWuVq0xzvc5Y8vD9KZ80kKlYJ7Am7roylboINey9DOGsUPbd2iK/48Rx9SVVN+
XQzkyNfISCmA9R8W5vX2oVfB7qDulgRV6NG9Lm2hYZ4bFZ3gxDBoItpx1ijplU0J8GAE3H5SbooZ
2Ey9C7YHeAnJCyPzFEyqXtXCkTeyR5Uve2wy14XZd3kPVMzMd+MTR5b7VdcqHTFrZTs0TPCMSXSn
bzLov0zG7dWSh9SzyK5pv8DmtLb09uSA750v88CthSrjuNOp1ZsrjltfQLN2HqqUTD/HDHxj0A+v
T/gBzFR4h5qtVw+t/Okl0DWKTjow8IcnsEldiI//SlOMKeEaxj2Cv+1buHscpDgap9nTBYpg7Vk3
LSRyu8cZkY/fLOfBDG2oDQS+K7+LA5JEyMRoaDZhz3/TWsXO22LdfF76tc1SRyWR2KHAleoDUgzc
ZcOO3b8/1yNxYZNXeJplpExYHcElnh4bZUBx2zxqV22jyhc3qZfPFrCl1uEEtu2jE0x9gKq17cxW
RLlO8oM4Rg3NOTO0XS0vXPHRxyq4oJIQ4XlhrUI/+6Am/u/U99sIBu3CJhOGTUgXK71Ttbx/Ujk1
Fd5dr6UyR0CphluvKYX8j+AmpJPtrqgJaQN+Wq9um30LCb36FZibdNDr6ASBqyVcLh+HcCLfnIof
5deVa1Of+s1h6VuWchpSsKuHV+1udUZKhLYh1d/mn2jl0SXyalAOqbiVA5T6gJU/8lNi9qgMlSEx
MQJmpYy3Qc7GsvtJfLv1e9iRm05DEoMYZMkaxrWA6xPGM6Z2UPlzeYaRmVFLuvtCsR2iaTdDHo3V
ZhA4v3ajROV++UzhosSjmU1H0Gx221BBQs0DbQiTT9LA7DbaNPy3zTruFN+UcSUz4EZK1VL8I5Dy
0cwm8YGzZUh5BjSectqC5nJkNePbtHBVvP2YDpHWvnAJePpcoKv5jhuO1f/bt7Z0ZIh2mjSFs4m/
YX2LXoBH8dx2oZw/9CdX4WCjxy4NKIvkX8AJSRKopfQsKmLNCZ2RN4hT9R/+JXeZTg7govdFIx8Z
fLgsjmxxiYxYw0/VhIVbTnuCFEQ+xol06sCnA10d/R05JRcWiqu2t7+C7uUcdzukvYYKdwUv75hU
O0CaO8HBMFw81KwHt4yANCvADF34nG1kCpSGu8tdqfEoakY8JE7N5nCYqn0LAj+OS/UimLQR86Bd
Cr5wxmNnVOg4MWqBdOBlZMu8gTUOi92f8zxmJYBKo/72JtylITyEESSqKZ8tSm5CjJXijY8PZjjB
L6oMIzV0BMEzckv/EBEcBYUgrXtQJxKqsyjIvyczieYocxbcZhGG1I45t5DII7WbP+JR/h7D3bs6
mivSEGowKWYfzt5C5tv6EXh+hirzSb/YtfdLjZyANyUQz78yfZmqCgpPQT0KJu6mT23RHQe2Zuag
auaxQ2D/cpNe2CLY0Obg6pZANCzKfMJl84agW2HceaN2BfNcNVudee/oTUomLQ8S6QSTtPxouaU9
LsvyqCfosZizZ/q2u8J4lwuKwm/TlYs2WXiWwlLGKhIaqoiNn5mQX0teYnj27rM1/05RsGX1DfsF
/2tdSCe6cPX3cVr0Pf9pHgyB0UIQVlVWqHdz2l5d//P0ZUKOZngBDl/fclGwP9rlQapF5fzouJev
T7dLopTlBcSX16bRY5xrgI2xQPbNbXjXjEVRGAGqgY+bCO8izA+1V8RSOss6mVRhtwMQN80sMszi
Z/sOvNW+DGfxhksBnZTCFQOtzVAZJunTwASQpHddWf4zG/ZWBzepmuIiROmQHqCFhOHukPEesLJ2
NZ6vf9Xv8tmqowAXJ3Ey6er1an8INpSgsUg3XKjxFnmjqAAO+uFrAqN/vVl641BWgzgl9kLWuO/+
SiYnq0U04wWoZN14IGWVpK8oREl/iNNtiX13yX08hDX9wrmtg8WoVHCG41qE77fALmXpuJFSwPn/
9dPWsT50x5WUP+jjeiXnKorZ2+7pJiV6M5WfZSarSmm3fQBYLfEL3wy+RKE1Veb+R+SVSsE2iNhs
nKN1jBgw5+m9RYDyzDDtx9gS4LFa91bxMAbh83G7x4uwaeWizTGZ6MQ4GUYTXqPyKbYB1v1mnVw7
KuLSTHQfiuYA7rpSN+h6/pPCkOACTOpwdzgBya/92ZIv5ZxBj0dhQmcCPIxR2WyZK4LH/uuiVAUZ
RflIi+a6W1o/e4uPJonnvfyt8+s1XDS1L+Kc7G3gSn+KegCL2624/VhbUDkqfdgaR21lEEHEp0+R
sTSUd0Os0ud3gNOZPbYGGdVyu867k2QVOUiHF2Z/DWnJLzkqaHkJXeoiAwzEWt981TctFA3zxRXe
Zx4gjN4LJafyzFJdbIS/e1uJVObeaYxSoxV8PXpBO0PAsO8S8zhEAptzLObckUNVjns2wAePxGZv
i25b+yDjxiJeUidOFlTestv+9oo+XeWoemUu2EayumWs0p/6sFj7rjh32RlXNzFuNCFhQTj58yQI
/HOfUQELhCbW0GTdChokH6pSdtMwtMa2Qp7nmtUiBVCM7v1aMjYKMBUWQ/8hybSaMYrv2McS/5ab
nWp7iNMYmVqGgDTWrnP5M32gZ5p5frAiTQudJ0sFfbz/9x4Wx85T/+8I8OJVBZdRgSZMOTgvM0wu
UmZEZM6Im8OG3KQ/5a59b7wNuqmgoaZqrbF/3bLIyh3pzLVkQ/qlExJqe5IzCr8ynLfIik7CGi2z
/nfa2sEGE7odyRzLz2nGO3AG6DIN3JPfMISVjFGcZx+gKVdiaGc3/YT28Qi0DGdJy8UyZrDA94Ky
9EPtbk9xpr/uwqlibHWnWZzQxPqBXKFmK0sntjaPiehIakdsbScdf1s/yyfyT+ZBe9Fy9+DHkljB
oV9+x6QCvyiK/s5GVhOLNRD9jG/uQyiuWCYsW6bZyjqE2JMC5eZ7/5O/WkXzrQbZPnOKT0XIHpL7
pprgAyaxLeFpWLs3BnKy/3m1eR4xXQFA2lZ8RiFj9TYYSdvi7Dsi+hCAuhbE8x1zAhrU5bHNRg2H
1cCF5Fkc7tbPOQ5K+69EB4DtEnzckjQz9guxxECkD2YFlUcazNIpHtA7/QLFEeB56AAiO+DViP5x
+YefEcBxz4vRcV1q9gXg3FkzKVhvKOmzf2vVlQvDGHpgkf6Didhz7DFN2VxzQ4Cz7f/8ZytSyoxj
pFundeETKC7oQynBnEI70n5cp+2jiRQFf7/tbVyFV9MajxNr2yIG8SFZiF4QqUUNvZjhocNnlf+m
dYT7kgJtrnr9Fk0UJsQsQ2vZaJ3oSXEzKWHpkzSCRUIuJ1iTp7wOaAwAQKxLtumjyWT5fkBy92ny
l+n11U+uMocaXirl2uG2jTTw0UWaxRfKqHGuR7QLlToNddU9pso1Sl1JVhR7Omwh8rZVgp7Qs2qG
HZv9gs14vtSK+oTJKuWdIbijzEsV8DanbjtVrm/gzxXJl0pTICr/0qvBIQ/kOeiRaaNp+TTfpGWP
wwFxm6YRNuudkjgZIOZO+Rd7g8mWn3ceqZYsjruBJloaSQCRLk0X2LsSmzddwfdOcX4kPMTPVfwJ
yfCM0cMyvIiAU+R5HhR97ZlTo84q4ki9Hn4QSA4Rd/zCQI9sGUyCGz0SdN+xRsvZcVFYqMzBpriu
kiC+3PmyI620zp5Y8vf6XWIjnqm8t5H7sB95IFVkDAckEqNNIg9WmYxju8BCLcPSyxAKnoJwT+nJ
RelvsDVR2J3EpNOZXsdKVtl7s41xuWKvO5ZJocilMGrLD8hTluqYrZGF4FZwSezjDWhEIfc+6vsz
0zHoBlEGzg0kTMu16f/ryGbw2zFVxtvD9YdbhwlYZswlW/wuhRtCSlxcsTTUOyJJzD/UreBYY59j
Rl4J7lpQBFnzDYT9NExZTr4MBhHt1zJC9Bjq4cikkaxWRZ/0Gs8lUWHbKBvV02l4Ig/i71cVruNv
yB9AvfPmG7OHp/euRDEW+V1p6ihS3ilhyf+NkqsJYbEUqdcy8qq0uLMs2zBjmVSNmN9W8m5AZW9y
jp9uoScBAJPZewyFBGlmW14lfVRknj2ku5lEUMHNwCtQc96LDqg7WGEQd3XkL7+vPHyWSZ50vyK/
njmP5ieBI3RUaDoQhrjQ3G6JWu5y88eufm+OW7t0wghZadk6OoymmPL/faPMimc/ZIzFP6r2eASz
RWsDLaYvEhHYymuxmPWXZTZuKudPqT3rlFezLu9zsq1oVUi5j7GYuCAaS2himmppr8V3wvMvk0Kv
fN0JjJzj1KE7otTcM5yP8n7RAvM6RGHKoTXWr0zVpbCRYsQmVnVvgpambOm9N3piqxymyZUS1kgi
usnP8GhoJ9Qrd1U+KEgDosuea6Al7J7bOmkjRVT4vPBABwYncO9eUzVmsZ/EvAVkrpkGDPHfSNrS
I84uCfTLmIrdXU8eaKJ+Ih6bvQByGkrT9tSO363ptSfv7V3M1qe3AmazyKtVPwbv7KBjSa6KHb7l
lXrAu39bTfSzzjBrzylRtsQaQrLMgh2jBnK6vCDBVwGJH8M3ya5CWzIcn+NwReLrXVv6WbXME5NZ
8zmGeAI3mvyY65xWR5BVwksKQP8vaP2X+hg0CPThlr6Z75O8JaMdvh6xv28s39FzDndOa9W+NNq6
XoQA7sDhO2n33r5gNe/7eTGjSR0TbW+kI3DZFSBgbLnFpE89dThbavpkjF2MsJbotWSZEfBv8TZn
3vXEeJpbgmOTrnHcc4pD7OaaBVmcbVM8e8l42vSdew/gK29qFHS+aZ3WB39fLyx9l2IfjmcwrsYk
TbN6ymxJ61RX9eTGT6+FIzuJKKe7m1gs2Mq0JBAcfMjh3h8zskWaPfdvYyTPwi3ZFaWaSWS7R+4Q
6EvxI0hm9Kqv2VJKFEEFBkKuZ8c8myFD5qBcBR19XP2LPcsvrA8sGVhdoeVRdXfH8mb1NwcQ/cda
Hdn7VQQqSpsPnkmqK08LfPekxRMOxmOW0NA1UCMK/+5n57yhKxILnJM7Q06S0WPT9tbVe0HJQw57
bqRE5pEa9ryAaX0SSYvPM0/4igxrU6jMVh2fih/5CLxim2TmdLD4sW5SgUho6rQx0swBFHfYjjZX
7HU6/89X0CylGcPdWTaaBEODhX3DlCm4x148hKrox+zNJ+z2IWP2PEGHBQvLpjq7I0d6XRYHXlSY
FAcJditfH4xBVcPPFksCslcaAJr5oaqDNS1VvDeJhC7yN2OtN6v+B88vWWjADbD/1o8W5YLLrVgx
JvWL70GyqsyPwhEHN3mpTKS/qeoTeuCzaZtzArzBSlue/m17oVmKAvVqUOpU+zC53PpdfgF7Zn7j
665n4mauhYPtZdkzvCahCJmihk7BQnlxi/zZV9ELaHYh5vPWOQxPUuB3WsMbIsYmk7tqH7eqzFUD
mqufYeeHrJjMpTsdawO5yXBv5SHWom3jyDXV8MC2CFECMoIo/M76IWfbCm64pxtPjuapSZ4xUWxk
6mV8J+9SK4lC73gkK35PiGF296BHctj2yynYQAtUiLFbDyJ/IAiEup5M/x4wqSB5zBeZMinbWtDI
7H3O9xh/EIoQdDIJ8+W9iZS+DaXU0qeba6XxMGB5uylbBzbIqJoeIeAibHbjOnKTPGuX6nFpSxWC
1naYByURHXeYo1r/aVj4VImLn1Cdf37bRBm2dWy7hJI2qu0L+F1K09LFtTNPa2LZIY6BvcY0IyeL
3p0v/ozoaRygd419DB/rdGT2zqmdrtlUdwE6zhX3ILORgea0kx7tAHErBJ/1TTgLF+7ONqCmAnLZ
yCNsbstwMPy3bL64An4avNTtB3zjJeXVOsk/u9lgq8AZg7tToSr9M0UhKJP0xChAzj5+ohsBA1Yo
eDPNAbvu1IitPsoefogf6Nzah7C6UkLnrqxTcVK3t9vr7cCvNjlzUMezuNcX2Ra73B7TPFSKX7Bi
VWRHGoYtObtWMDTvLQK2X71xyKRmnb0jkWAvybNs1mVi3LNLVqYv9tu4+XMHQraWE6gRYG85WzjZ
dCmMcPJiSgQqgsUzKlOJHC6jEILuRq2BqUhFBr/M5A96sc3TvSFqnQ9J0oDpNESXLLgmR01HhVmo
+kW8deOM92nNxHhcQ65JutNWrkp8sL3J+PfdUyVDOew9l0y/ypaeA8RCdLnDaFDCD82XJ20dNBMt
lPF+XLAgSu74nT3jPZwjFwqjXq88wmmcoKhtdF0PVYyoQE6FREOfxrZW9v8karHFzG8TT2naFeM/
ppiMJR72XmhrySGIgW6kazW+2UojEzMsWzNzBrMlqyZMrTz66Y6iKdRnbRXEIKFkZjkaaTPST5nE
xmmIV6ynAvUf0JP4Xlq02WIc0OWSFEBaTlyLf3IWW5Yclod5LcGbPbM2NvZSP1NERc3amqSWmxpN
yFfXxg9rBLzkdlPqePe3h82JszmuMW0hsnbjIlOz2YNTA8h8VcXnQNbrSgRE0HhibgeGD/q+KPcQ
yJNufBzTCOoGEcvWxAspdLd2BMYgRSHTMzQgqg2qfVFmAhihHEiJR1fuSpb/wtg4NTsvaQscccEA
uGTDwB+CnYqksChGSxRlz6UKh3W9bWlnBtVLmkGJjMkWXx/Yc5BMKQKBuV31HcSVJUoNyfpyWL7K
+2pVTdVeWA6DXndghc7oEPP4lej88YjnSupS+mwMDgxUAKQ27PmSj7YSYj3B0UMN0aoTxYvS1w/m
lYrtG4uz6sAHj5hoDJphNkuxk19yqDCUnPTr+1I8ebrUTEaJ+i0yvv4IyhJXkPccWIyVwB30CXKF
IZdvhV8/HoZyaLWm5gDUVlgEukw+eD0kahR1vkerqhLrHIP/xbKVn1iuGx5LsdQjRHfxo4ihl9aI
FwGGxU5aRbJ7ZG8/NKxvyxSCnYPakTqIYH8ElQ4TUX5BEYWMBitFz6w0msbQhHnq8eniDkDE3TW8
N4A1ZJw3Z6uG1wbWEGCVdYZlYK1fEqhPz08v3kn2ffpn6R3p3mPXhqc0XC4xt5MKLqv+9ELiwVPM
1rom5czJWvhbre0tNrtlmq3KArFSC6QCyZqP1O3yiBoqvVWr1+WplsfujiRIRMnEe/Wxq+cwFVkl
c6xdmcj9aJ+mqQWEsTrKcTPgMC3qtUDpAwWrYPld97faVqZwPIFoq9JctIGvfxzD4AJ49w68EIU9
UXCqJZeVYLq/wUCg8vn5ogPrQHOefz0bfetPF+RDoh9w4vpUU7m+i2z8qhuaY+I5bEi5mofBiDW7
VhChOGUqx8BrudeVDwKtfwUNwS5XeDidFitFDWFFNa8kdWydd4TRC0fcCJ+p821Gca/VXWb5ispW
4AGp0AllPIPphfWA/vCeEi6x6CevDF3aMQnN8Gs9MPXx7WVcvU22RcPh7l4SqlyEtKV+5fHF8zJP
pjcNqJ+P91V9PxnVGF3oAEGxdcYvCRi0rWF34MOedLpHuNMeH9HYY6QpXnRpWPUvbykfW/SmYon/
1TXvi8GJblKA49MyWfmDhjgV3fNEijvrlfhZSimHzxTHQGAwm+vlngZeMNMyNvoheK1aNztDKLXm
GfGsk0fMZMUdScINiNj0b1fxKcb4XrSwsERAsyTIihfSLtj8VggPmnUVdIjBfZSu0A6l3DqunBnj
MiJMiHA07s+TcgDf5DHUV5FVh8riuGc6p28xyUf1D6y69xV/DpHcUmlURubvYoOw0vTqWzKQSDaJ
DY047vxqt3AuZfU9xjWkfPuC+djvgOk02BCpWkiD+fvoaRQ3a0R1O3UtLtHmgy0RTah6Sw+MVCOF
xBwljXa1ahh6GxzcUAiN8ON7dPHeBfl7NhSm+1mg+VU8xgt5udXbO07HflzuQNwdaLSytnYCPb+N
LifXCFd2bR14XugLcCfUy4k/h18iX0CqVA+2enGjmEaLxCNpzDiO26XcUTT8G6KYpy0dGF1Evd1m
6vXeYXSH2r+mLWYHKhCXHud7GCvylroxhtStiEdaFdUWujZBL5R/ZgAoKywm3akiGM3J+nxeRnyE
38ZkyT0DZ1Cp6NMo9MP9qA6GeH2xeG7V79ruUVhX6I9K+5wYtrdTHam/b/ENBvln95XVxIeFAtD/
JcYPir3EY5Jmf7z7voIrLi/xD/mUeZkZ04/irg5cFU//rkvCBDiXTXBfz2rQWFF5P511wEF2LJfR
/Waz7JV9OAKp/OOyyCQFC/27J6v3V19vBw+K0Q/qsEFaRaM4rAGID0i7SgG4MXkXV4msVcGwxUdL
XJoHCluc8EC4ipQp1XZBCJhLAuDngETE2di33MJcNoKQmCEbQ9yx4gPl0J/Y6L5ZSy85PprHF+aN
P9eNT1bPo+bqqK2AqKMw0IqaTiNwlThLyOrXJjHhdroHn9iOcMCPbYQpRvriM/yTRKBDgbmMuU/k
kTf2YPq9F8KxhpHFrAh4Fz3oNBzCp8WHnW6yE3KJ7zwVjb407ZfiMSCwOkVbl14IEGRtOIiD0qiZ
3VNrVsvCqazAJmkvnMqil4leY0wSLaJG5LZhCWlq62ncGAeGMLjSqfw5TPCLZHOpteA8JRhKUcrT
5LmKRsH43Us1eV6uuh6ZMiM95OnJu8B2rUeIsf7sM79D1O03Us0308eC1rXlZvgrshwDtw25/Pr6
eWo4BtwOqwIOO0Plbl62X9hqKXNdguT+90pR5Vz+zTPmqIM3kh9p0z4Xr0R1EauOsF4lRy+C9zUd
P/JBv3EDE7Oa9wsSxdbtjkscjrafBdKwrGxJ8xz9c34XTAwvfv3EsnAjGV2TX5CNh2u7X6msile7
v3MTFmMSx/rWlXGVAyrytkqTsQFGYt3JWEzxXRtkXHd8RBD4qI9vWceiU515df9wEsREwaEDWlW2
e0n/raQbEDP565fbprghJx/PTMsR79zQsyS0H8RyXhdKl2GNHZprWjJ4YVlzodb2iXE05bHavPAy
OerKDmmO5crt1L0et96PHFTH61mkNo+QIDYKcV8RJaVvs3qIhWL+vmy14W3R2vILodvCK1xvEp2P
JpmPwCZWSh5C/Un9eowHDg064zQKRgG/CqeobRxcApx/r3DOHHGJqQj4Bok5BiF97+TWq734BLP/
6WRWQKM5Qghrr9VOmX5zOoaJXqYw1StnjaXPa6X4FfI7+bGLMj8PoiVkTyPSVoyUF96TJ7zyu2Hj
3ctpnWZIn6tGQDujA8Wdd/7hG9aFwfyGOdUfcKKuEDjRL7cSkZLNT322Qq/gc+Car4gmIdEaXNVI
wRwUk9XGkNQP4fOc1ombUeHPlxzqbl0lwHGrD8M14h5AnFTbMhxAxPSHc6vlsxW2XIfssU3ZKNwg
WrTt4wJqSuzJLYreH95+my+K/FNza7mhM67wsCJVMXZDvb7DuCLo8Wn0BZYyXevKU7JwjEYtB6AG
UHZoC4y+ylLWDd+4L9vAwZt5j6L3F9otudovInmST4C1yCUBMaV5FTQW4bHIOVu/fTiCxHtus+lN
85aSXMbBXMh+QK3UHzzFoY6B6/QtxCR6fTFxawhGKr9kc9DHcfwtPi/QgEdJDP2tNLmir9TV+fKA
DQmKX78lnr277jbatAFvhDG9H24j2Ak5QZs4X583ogfereUiBw0gclRZpGpS7ut4AkFYmNpH5rbk
Dp8HIJeoNxLS+CcN+JCwTn2GDKZtQkTcsvzPuGoIhqKIMJ/oT5+UPYh3ofnr/jHI1BmZb+HFNSPe
mjPGkdk+JLLhQe6JY2mC/01/KP0G6hMjPqzJkdXA13gJddsy88erRVhbQ0a8Y1pxUv98+/AKXrcE
D39ORivybYJ7qKqE4JJuu2IxQnftIi33J7QKJe2nmMzz7mcUCVSV+yBNK+e9rsCiVVA62JeX2FIO
+SOUpUmitzoXNl45DCkAYHSgoYMq6rCH5yQDNbW4hysVSuNKfIRgn/jQhdXAALybaDB2AWmCHsfl
38a2agc5lXXuVrE5airhWYPZaoi8XLm+cST9ZuoGtV1boH0CWMBP0rtvgzB8ZKBgjydN6p9xR4sh
ohmR8BnQnW3UD54NjrQmrChiigaYBV13g0EAH5HKqfnN4K/4vymHtSdeGuqc2GNWP5ie2zgw9jnG
PLSbUT8OyCmmd8zMAgHR4cZ3COmhUXWmDjNGIh6nTG9BKVP/8l6qL4/8+ULVIZ8nId8RPTpKlPJG
tY4lelKFUpnZlLcoLgRsP4VWSlCFxwMzih0hjrAqIniN0DOCOOvAtm7/byFuyevxO2saPYQq7QnI
1TU/g5MwE2F7oZAQuoVaQ88A7UxEoTS0RBMdgmLHwzph5dR7wRBN32PY2fJbWICUc9MyWqF4yXlC
G0tHHxtmvIHZKhfxS//VFbrLq2Czh25Rb32/3FZAzfv2ZMppMa+aQR3ScT7G7IuFJMsF0NcAdlvQ
4mfMigLAL4eMVVnUvU8X6SZCDqAPDvT4RPdZykElp6FkcuyS602Khms2E3Ud0+5EkJSM0LA3jtKp
mQF0/wYjygUxcm52Ws+CELwRbZSJqikkgihvpfPnji7l0GZZiQmuxnl8NAzxvqoh2QjyZ7n0QdeQ
B04OIuRp+3hOhOKrxaLN2UK1eGwmRFomUAUWDrtFyGyq/P5BcsUWhu6jGfrdvv50QTFQASWPPZ34
1lZdWz1/UUdPiSp0a73KXt7vFJ/qKTYj0qEBqSXiRNqZlIZhOPog42BhXijyNRP/6IQFPkUnLsl5
hmh/P6GHbk79jK5LHAVgvz+4Ch0sRBCcS4z799F1VJZhHmW/JvpPXoEsmvTJ+mrFXPLkTkuOtGj9
xwPI0Hr39GpeJ9rp7wKXYVkdNnlFqFG+k5+sBx0xg3dTvCP2UIeL+dmpW/7LL449Cwu+SG3CxVuT
SN6K2stY1ZwtHR9PJ0Sn6GF0PIm30mEBkPxt90pjwSXye0Ijk6ojskz0tTNZiXUVi+YLoKbniuKv
Y602yFRuM+F3Can7zZa8C3My/Dx31wOxn00Dx+4uZ7WpdvrkQhh2chI2bj03/zqMIo+42cqqyBr8
HkVNf3riZ5/+WiH6fEutoIKDNjkzXkz0/moUXcEt00D65eKifm1L+B4hyfnQjPAG9oHlS4Mb2+Mh
SeENZeHMI4sQz+kknTEUVT4O43yVNf0RU8iH7UVCxCRFpkFgpBteoV9NqzGyphz+F5d8OVnJDgm5
R2sBreWs+sjneqTO2FXeqnB34SsJoJw7thuP7XvCwr+0bm/pcvoALeVVsZFIqYcn75F3DcB93GhK
sUbVqlYfUDToQgxgJl2QZybzlWR6EhwgCbUeSLUe5zmncKpdv3feAoP//PHC4FOWlatwX6WAdISn
waTOe56OYq3iIHn3Fa1XD3CkSQwUnoZ+IvtIX4PmqCJIeNqEJ0eRRgKuqBUKkUlb1Nk45cK7j3Tu
h42Jg3VmnLsFFKm32JyBiBuJLCg1UbS1pbeJsQzMNwi3arfBi5jhzg8umOGhEU+3aPOt2k7TF7ze
wq5RrwfOkgi/8YOdIBoKcxgbOcUhTKqE2Mqa55AMTRB02PF0/pjlEsUZdbM2rz7tt6DVMMgiO+I7
PUCCV6asSHrmTbaQ/B3I4sfUXnVRpJUkCnvt6s60HYAyQ4UHvblARY7mMKIHHYTnjQHIYZoWrmGy
mLxyquRo+i66gqkD/Dbqw551cOzCTRQRI5ViTzKVRDUIl7KaYwyu7QV15gyYFHETSObixEHn3Rac
G/ThvN4rNPkB9JBtQXwpRyHeYAfqLDVQRn6Ua1bFd1HXoxubBCRQkMhxUeV19NzVkvOrosrbvwR3
fwLbPkiv2+pSeb64K/9hrNTRIBcp80IDZtVHUwsQzlHH98f/Ymr1veRwbXCZmlv59IG7I0y8bYCe
gudkZh48Yb7x7eeqbD/aQRydK0hOBvxbIJC0z90Zj2R6l/37WBxWZHzbCcnEdaZHunndQgVW+Zii
ZuOkO++o0aSa77X59E/PysaxLXJ6urhtVm7OnLoknkHimXqm5FMlseKLYNF4QXJCyXmyG5lltzE/
DPZJULBwXCqKcA1jL1manjLIwMF9xzpuxu7PL8NbcHDNYcRSGW0tghQl4CJ2fD0Z8zahhs8sGUTw
Lmf678Wv+qNb5V5/vFSNe3i3KPstjEI1ulYPG6+WfQWuyPc8nxmHVA973P7K7Zp4Rh1bylprAWo6
JKEklENdrwyCda/KGYmY3i4MrGSQYl9brC/ELK9H0obGLZ/65coL/qHAiK85YlbpRiGeH1e8pmpV
OdUmMfsxBo1QJSrqmspvtQeHz0YG6pBce7gioInFkD/0lM7POfldcydIF2lqY3vzANYv6mQZLq3r
YjCBljyIO0skwyEjiqB7w7+fDHASTuw28qPTEdxy/tuKoZ6PKbQF5sfuhOY8J3eQ7QtNJNyVCC/3
6TPbxarX59pHbIAteRmzd6Z+c2wJZFCQpwtnhZazs3ftF0m6rTwSF85+33xe8lK8Jcnih+7pI3py
hXbdqycqtcbBRBZBtoeSsxkvQxLjaNZBmWVNNo0YAuwW1ts68c4YyAWwfAFfQatyZfVZAY5TTEvE
PPdSMhW29rpwr3r8lQqyTOZaKFcrocEpW4LfJmB7JEyOcdGAw/5oyGl1jFteWQFkm0Kji+Qfr7We
Wm2sSTQ1cljRDEK7Ie4ZmjDVjC39wQF5KhlvZ6//gixRAqvGDlLJ+cefXocwlHENicvMIFCT4Rk+
e21FYZo1s4AT4hexojvxPhH7Ad3gXeHMSK3A1aoDscXtPbNHV2LuuFOprnJ3I0cMG3jC9WJvqGXR
5QQhWNpALER6+AMXoNE2K0uHKgxFrWF0E0WhF/Upir8C9a2Zy4DXFLKQuRqpYVZtvdhYdIfqAe5w
bmgZUVuiamtAsDfygNRqfWOOVZPHFCM8anxDqsgK2uDEabwQgIL9eo1LRxdmHn4hAtDqUQ5F6UBr
BR5vQJt8UUWXDrr31MqQEOUILg4MTXxJPxCn+ke3UEN8P45z925tjdOlO7NV5pYb89Td9IwYSjuH
9VogrGiQUlpxMHqslGpex5XbshL3p5CydXHcdpFSukL1koMz+LNYAFuAB+fvOJRgnqT2a9O8qqGf
Z26Kmp1AM2y0jatiw4lo/KiJDLQIOzmj8hSIh9bGwSXBp0ybd3U1ZycG48GufLB8kDHt+32lfqTO
dNb/x5lHdz2Y+tdIqYdiuZiYnF69BNSFenQpGPsMbQir/CaAn2SW/piyHRxWWWam/jVN9o3xqPGf
CjwdoZSn01spsvXKwdizKbyMicR4HlfZDckgNjPmIeA2Y6nkfifoj+4EcCXQN4JQqP3ff8RG1X9I
joUPs9Zo0P6y6AN+wjYRhLdn7uh10ssQiGOsLL8tV3OniFa8h84Rh+6OgltG6De3eIWMbv61leN7
/Hn/4FGZ0hD2b/P2gPJvsg+1rYEZQbL6PF4T/RmguFev8GA0NxsxzeJ/kBneSLbn3bVrTKmg7b0G
PtGvtXEWj0ca+Vp8VBImngevKZylD/MN5w+/mEWUxJg65to/7DYvwk+QTOfImfwZ5m0NK7zMmc1K
VPKrX45yFrsGEkm6pnIgDSpANxqTdHFIEoNcLgZMgQ9/qIdi5wXG1E4lvtpDvbpe23WLl2zV9fxz
uelnKE8lRkes/G39CRV3N9MlIhbhgfqXvAMn3aN/DZgA1ggaaSkRHhA2W/svC9BJVBbAfTkETM5q
k8G7vOMzrzfRQGGm4ZUCWpKscmdHl2AwP7apC4Dmb1pDcDcMT1miu8mkw/AenV9ljVWi8iR1dOzv
kSCAXliHN1iTLyFdiwlh3ieP2ZoUDGYOHMfZKRdcuJ0xamGkEZSRwJf7fXJvbyCnM5truJGPtpoo
gEAMUbDoLRmIx4PMRqIc+eqDTRaXVigtc2I7/z0SylTKNILEc/5ClJ5uKrpQUVcGNcgIp54s/JLr
sQdbKmlQHhM4J0i5M07vxEMTbsrqEsnoh1f/oe2tBThgzHsnDtqpdUh5QhN2ikPcjHE9vj5A1cjT
BQw4h67HzptenDTYa8nUQS89R5k0+cU3m7Xadr8lKEd/5S2oTtJgAONI1OljNnUlx/HrPmfcr2EB
jdKLlNH0xPIocGS4Q/X6HrGMA+0regeHO8TcBiH1YqBfh2Is2SqpFRoZoesMpFoPxZxqt3aZULDs
ZCGRaYK+hnqPdAPgmMwZ1AdAs6a5j2uUnqN5WPNxgvDWhu1S6ghtG0elhAGjlapd6YgUjGXXv6CJ
VwURllC2sUnrtnRdOJIAq1q5S5ToWvDc9ax1EXNI9VSPKxWCNYpv+m+T5Nl4Cc1i0EDlI1Zd7FoM
keLbLvLEzMUWEI3DaK8awxs9TZClclgH45+harMsBfgWFL41SHbD5WrGKOn9KbspLIZmdRZzAzTx
3MmAcn9esKvv/fjH4znybznX9nEe3m6SRu3azpqMB+RCpkZLdvLE/8P//lOcdWFLnRgutstD6jhk
2VLZF/TRd6kNww9K7ERFv9BgS/JjcAPw5CnKCW2OweNvZE6EH9+7RadLWalvm6gOEO7YhrlI6IJr
sDFwqtpcXtR7LLsdnk03dV/YS5xdpVqCHQyVWwtiOoN9Gzr+65WcsCpNC0bkt96rf8fR7p4gDmbZ
4/bhckTSDeBzQlYxWsSIo/JCt5reU6Bd+0XpGWsW4zCxClLlH85Ote0pP+DnLlJUJSCColbVdh8o
yvRe+En/Md7kbjR1vjlA9BQeM39W8hhckIlWv1DDL7vLSzgphj3zqe0WrLGKEF4U8sxrDpp3L559
zDHFSDnU0Xgt0FzP7apNNuR27YuiHufoRDrfFC5IOhG1PDr9Tq4etXQ7JgSzgTUcz08/eA59yUXW
YXvMXnx91c6oP6v52MBzmnx5uRISu57LzLDWKb5UhaFCTReTNDIlavVT5Yj/HDO8MaZKIGhqHRNF
7VYwSxVHWpk13Bv051VhgbqiQoSBCTMqkafzXVjn/XLFfSFocHGNxyNrbFac5655N6AsmE6Snud/
WWWfj61yUpsMamx88Z8lR8CKqdEHoLLGgkqdmiSbImfBNmybXOLC61TXMnnkREdL6pLUvO9kCcHE
qDMGyz3PeKym8LSyZPMyqn04NcUN+h/zdfTbL3kwV9kgQ6Ig2yCC+Qa6r2meS0CNvrttZo9qyYGv
qMXrvtdaYG9egnSQFz95s+DUEP6/aQiakz1GRjAi89qMKL49ZxJp4hPdN18maz+abu2EcP6Fs7+r
meKgvYIYR4chBGBxRHHKnC12UIlTFRGnFYxxPgmMm6lLprzB97WTgD1tcSrPjRCgdrlKxUlvmd5q
9mkwpQyk19GdDtg7r7S1FSUNrY5mpwgUI4UuELJIBH48aX50RNh5JhLru08tHzbx2BmYy3SR8ZfV
XRKGgSdiZMy8KGo4lzXr1YjkEg+x1IK7CLz8Oy9IA7d13xYjZOJ+PZxgiHHRY8sgpdEUDnr3qGbn
TS39G56TI2+JCxBl7eD7VfA1h7bRiKazKa56IJDd33mP3hFSAWgaHAMmh3yJdEMLdbV65WPZCiJ1
aQJ2xqpD8hE8LTuNaQDdy7OGHDguFEad7uEf8AUB/2UXiADZDWw0BtFsUjdp1OFv9R89DixwfVvs
Oa33kv4CcbFof/Z3YIrgceXWcORv922fd6y0Rd/kmZPou+N5LSlFhNvAh6HxAWjAVt/akjTag/bT
6aNcgC7dK2pK5aSEl75R40rNoaQp04M0Y22NF8XFgD9gmfg2UtOcScTCrxZ/2Ci7uHxUWpattFXk
L6MDyfUpLXVOcXI1PxPLuStx548NAeCs1gT5q6yQFWFeZ0GmOrBm/hPrWLJEi2ZEgpA+q43y3mYV
ioKU73Y6yg6KEOILQVW9HVAGFvi0UrXR+GVEMq8VMT7Sdys3z40ba77iw9H1+3eFPepcc/bYr0Nc
BzLphxNlyWbZR5F+UjfcRooUdi/3WgKnj+9KJCbpUavrv72bnfFG61gAJz5FncXuQCY7web9uweX
6wqiEroJDVITwYkIMkPgXclPV9MbvJ/IR1DBs1mVee5ZIzTTp7n5qfWVPpulJIV3ZijaG27VOXZa
/QJCS3deFFvRu5GzlGhn+ixPWgk74RMdvmYzdqZrc13WgusIVOESAKo7zc/Z6+tE1tgjWsX27boL
gRNOXtOHMouyfPTgeKBNDFfjqiUBXs5Vj1caFj+ZtOhQUOzpRR2p66g4TGVaEmKsWy/viCzpMNRc
gsn8hvMmjAMb/k4fTcfPaH2hBDKQ0hkFT/GNniWAw33rRKxXBZHYvhHsP7HqtP2JEh6xv2+yPX0S
yrwS35lty16YoEujEIMTd18pf2k9CRUBDBkHSXmSzlw7htjxhLIR2FdAvyA4fzxz6Leq5mFxYv13
DuHRON0Pw3nT0hzTFncfaIftWLo0DuxYG5Or/39RWMIF10Um/KD7zbCuJYz56LoV4F5AjbbY1cKF
7XH4W2jXWF1mVw748TGMXGSFWFuBWn4or71pAPY1DU6wu4gPflykkQ7OUCqNmCbnjXBcj0OxfUwi
WnCETkiU81aoC+svMfOmsQbBqodoVJV3HNYdYaIqlC63ZzG4PYQaEVXJQg4kj1o08Bs2/QKfQ/vn
AqcgTkvGhR2ex09kOtwzepUXBkZ3ix61bkm8a9zJxic6kOKpZWSkEFk+OPcpahLtC5tq9fGPOc18
Uaf/Cwsp7m04ZjChLacEWvohdpQ/mSYCaWFSdWOe8J72CE7G+Py8vTKRwsXQD3DXDV3yaXdwW6UM
a2lK3xp/DYDrhO/JwA3tbvY2jkVZ/vifXRkPRz7/+leK1VlSXF1OKBGSdq0Qjn3jAToHOvL1Z4Pi
PVppGFof7pwhPp1g21wcmY0pkQ/f7jWg66IxsyMl+S4kKQbdElNX7ggK1iDSK/ERG9U+pbbCMfCY
8knY0QGzmipHH/HomJnHsWJ7Z7dJXyMy1Hb9i587mV3Vx7OhiLlKWKEeryA9h25yYPdO0Zckr3LE
3E1pM44wtpaM6ZAKTVm231pKg8J436oP608onWfnme5MB3n+DhDVmt9dx/Tq8bAViOCs8Fl9muQN
zHdgzC53DlUJlx1UcA/UHCGb20Od1ROfNL5nU0vgGZ+ZvRA05Ppq+7LtaO288ySFjQZEMqRP5OPs
p9nhI3SurUUqihCAap7KGNgFYi1NRBVs16bu8BgUIt404YOSMsEwl841zR0g16sJI8tDOSShVmPx
GCxVNuqJ0zUd2cEo3h/LdpJWz+/wy+7CeJGPEc5eAbwjfnXJ2cCkEllGJKDGvBzm+ucfrDIOkKS2
LMaXkwGWGg+UttQZJiCaUx5jl7pNRltBYEO8qOxv3JdN4fOh8QqslsaZ4DDM9YxOUYyXw2amuCio
yIBpQQqjDQtqER3a2wX61C4l0Uko87EcpK5rwEXv9Bj3Nk3+a6H8Erpt477fEL83MXqkL0Amjr43
QPopYPwcGNqLsZODSlC+KuY2QBl2rnSJsbIBWPVbIKVHqyVbaw3AYKGJhUMaDL7ehSsKo/5k6m5z
nctl3zixHp8QKmp1zsxQtBPHJYnZNr+hoSCPHHyM6h5LXM18LSS07QrH4fXBqzw+mh+Xf8Xw2q5E
TKGG8SRtWSmVkigDSGfdLjHLIgmC8rRqWEP6Ybh/WHm59aRVLZU4ltN161p1cWo0WzGnd6QsjqqR
6Nz/TStAM9k4H7/3CtOx/0gVuXfMly2Z2bXuWFzWX2gn8tBDWSm2lXBoCP6xyszdTky4llRFbdc0
XLtqBYuXhohDMTQ6PXb9wc31p8s1fQHx2s6OWdNRA+Yb5/DeHZjqz3Y89hM44JwKougYL3D7vkOR
8gnalFJjiZvLA1mGpoWdxg1C0Ngkx8zYq54Ee9j+gfL+MRkKuWwLg1uaVVkN7Xlejb2djY75U+qb
xvpnuEmebVb1I2QrCl97C1qvy2FvngVDi2quZCVfjovqBc90VqpxszZUyB+EARb8gX/drRn7FnhD
vKr0JRF4MTqTKH6Ud7TKy/mmS5HRoFZ9li2DeVJbafcLHkNTEhubdNNOpwlulcRKksM4evLxgwN0
3cez8gmN2TaEk7CTeLr2bsxc67hqb6n0YB++junNF7vQpRQB7j6JULXUV8zxqBQqJSxEhyjF3XFh
TTVG3DTGve/O+kz8QrxqrMBZufFNLPG1O4YByOlYCgQH229AsoG7SFuz3pw+WcAMz0s36R72gP70
cjARKXvPgQ/SmaeNzxWQWUcjfQjOZhte1zQfL2/KzF7FEvnnZ404CAAJTW/9EsVVB7oItpnHV9jr
hT/OdH/L/XXPXNqjvOHtVxJyM/hGK4apRj2bHnp5K/i5QGQamSfXja65ES1BYkRl7emBV1Ou9Qcx
AlNJlbK3EMyy3q657kp/ufqcllX5FAeqG1r82mPcZfLlqKkFPy4NK3dCUhymQ57brB6if06Yn+/G
BvKUiIM6gcwQVdzeF7/2mNrovPLPtn+R9YJT+YArMGZt4AaYQiPXgi0wFUVZkA0SBeQ6J+DhDVt/
abFDNiRlP/XNnyJPJ/9PaOwiOnq4RkLdrqGJRZnet1fF9DRSfymK4UVb99GdM7CEXakNsvkIX7fw
sfTnDV6X6X+7WIPqghp5Hp9MrwtNzZwKUetoJ5+d+5XhbPLEV9ZiVwygdIPZ/n53er1KYNQ2ASZS
qzDZpnx7WPyxkAPgU11UW46IcHx2ox5F3iOxgCdpq91pEtBx46/jqKsdTF+cYghQAi+LFkj1fj7t
8YPAW0ZFMf77uE1CHjIunSH/QOkcPLAivFQHjAVrUI5WLBZCEhnI6f7b06MM5C3l+OP7hvw3qrHY
45XEz/N3YO7lGdKIcAT9cv/nkBzKxgnW5excbipBrEjCoTy0QQ4/wEJwwKW74S1b8mmJpN9XxtKK
Aj/KwY7hpOES0f6JS3yVi05Tt48PynNGLa8Wtz/I6SctBwp0aodAuiS7zIMA1KHIwgcM+dz5H5eW
efiQQTkzHMRRVlBjab7F1AxWVJUWEW0v7yRxL3cSjNqKDzz9Ybj6E14576tCvSkBeoDSBzgLahQC
6sAclvJPsZ32cjYjszEw6+9q1xGD/4Pa6AWa7Jea8+FT91Re44CFKYIyy5BUPe6wkvEsi0TerMmg
0n89MG7uR31ZUzrBQebfNatw9/TsuEAdb5Wl7ZFiqCts4/wx5nSAF7nnS7o5AOWL/aqYKCJ06fyC
V8/82NuDAXkEuBrWiuRRwV4OTpXDm++BjvCVeVrGL32pA2fI1lFEJjKdt5iaZVeiCiYCNNk3S/8o
qy7LjmAY2YzRNPp34dfwd8t+YkENCF5jBYkpb7oOdhVxVdnrTxP4tNdseTgYMkl3t5zxyFv3wnxi
1yM6eO8oauGPXgkdqkFkXDnfg6HfKgQ/QJmgKH3X4ASEKSDuRYkb5Vd1/ms1IaNX/WEi54a6F6Ti
s565S0crCB2eXE9NwARgdeVAf3DQ1HrbslOA6YhpcANZbWzWisC2Pfkhbppxrpuqj79v86l/ymqL
0psq/iVBQ7YM1PPOeu0k+OoXT4gMzR0nBajfoyqQuHYUUTF3dHNvXHFubZYmr0jaVOdWz5eBseOT
VruuZzlYMoa7NmZSfhRoYrK2ph6mqS6P9UJaHvaGL2DNbFx5TgJLqQGKguMOrWBBEJooEpL2J/zA
ti2zunZQHSEBUzdhiusre8M0ISSANYIqgvqgw/W2Aifr3Lk076zvvB1mLqhLsFWk1pmR1v72B7uQ
jpyY8pw2YVkck3Z7hgF1Z7VtGzHYe5ASu5StNHqRP0HGGhDeDutfCfOVhQQHFZXRgudOOrrafWIR
sD2UlFnD2ikrSfvfXMm+I0T0nienN4Tthsk90cc+eH1j7mEVoK/H+b3LU64Q7NgR7anJlbNyaK2Y
LLrVTC4flRX+opukHV1pt5AQejn1lvwzuTP0nThe6z8O9jyZjU1RuSbPkN1Ul4ov1NnvGIbP38gu
wwdNlvhQjos9OoMBUYPzjAXCAGNXoRT9j4gl5rH+8GCPh+9xYY0W8QlvQfN2pdK9wV6dmJLYXHoi
vo/1SWbBI4VUgMRXIsxXshwHHrQ0qWg5cllisi3w0Pf5DavXRzpOVsZ/WwvkMAmDHMNxxLVWO0pA
5GpZx4E8oAfg+JeEIDG8y6KCaooftubVGGpd3SqqnxyBP2uDKdQ+0OSAu62oQUI6dy9kY4NBlsYC
aMiBelQ0//8du0s7oHqFDnl2dyL612zsEGcZ5mE4xd3JQmAya8MWbglVQ0q7JCev3QHc8eE+ALrZ
QSQS7sdmgmNZjy+W1L9pFN1Uwfz8YZwBC9/oZ0ZqHL4VnnasfR+ssKLXRtlvH4NVta3qpNyWlejd
NaGUsqSMkafIF3P/Cpb0VbDGKVuVYebGo1xKD/eOjbGioarQuAC+bJnbge7JUbs2kRUKlOJsVZFi
BTWzFHQEhOCUl1wD0dtNRV2/14ahtx2kwSv5pAExCw53o1CRENGf0lNPhwjG2dz90gUPaPIgRJ4b
vuGEIHZMMhrQocN406BviDmrZkOEoiPdAa6BYy43FFuvyAK1RexCJCydheQLiromGQHtxL0XQFl1
gf9Eoone8d/ZeGS7gKEX0JilAqfo7hZQ7bt73jbpXRzV4309sbHSF7vQNcK5jG3+x4swd8mUzGyW
y8iLr5SeRRiwVBTiR6FHz45BCU55jZO2mXS08EJBAucy3C30qHAi2lx5W8yxlsoUH3IR74L5Dl3u
F9V3aETuwq7mzDnAtxRS4qO0kD1VH4eChv4l6Noy725mA0KVxJOsPoIaf6GXbWQNv+aMp/NMvdCn
2FCcbJRt9DMGH19UuQP0jJvj5v+RfDptgtMWgCM3+NYq944E6RlL9714qEsR9TO4M9j5RwlPhMuP
bXt/k9/H9O+49LeW5J/6roWfQl8kDdjQHSy2wDYQY+DgcGl7UksT1aW5miyrkdYevXz4P1o09IOo
pRlTv2F07UtbJXAPJeDuYHeVLGkTsv49xxIiM8mCmSj+DBGtqp+dLNpRVypttL92lBC+WCD5CGTA
oHl8T0IXUQlFnPJrcQZxOolFtzxZkte88THeR/QRJSogYRgLDzRp1JLdki0nXl83XaQMqb+rZh7Z
cJmds3CtKevL7+dxMHHbCQZeDD8CZXECEhlexp0b3P/Cm/xpqrbbxVnTVit+vKTacSFT5NnH2ksr
k/+gqqe+d8IRVSS2guqFA/hARWghcBjOoC13UChfX+AIsIK9DwbiWuq4xEXgAcUxVx6Q0R20/Ohw
8CCqwVkps8yl3KlFkh3frn39AKrtnwU7aXWFffi3ki+UKbqXC/EQUQd0uppotqhN1k4butMDRxhz
mC9GAKoN8K0db82nH1Xb/7XmgxYSvYoZBIeoScSRaRr+rcU+EfVX36W1DgczyiRJ/v7Uco2rrISa
NDMwQ0w0TP1hiGO8pP/qyFT1fLTs60OPaw4qLVKdAtg+AlT3QTWn076siObqSu4cIZ+oqSjTvfz/
PFW7UVKaTJpRyEXvxFvGuFuvlmToPF93FHhx3FmLavmjon/YW9pCVWCghHX6SZJnyo5oh62s8hrT
3ZhCeOnJQTACBLHFUMs9J+VSYAKKd3JAg/DCVUUWi/DNzVP0D0NraZiz18bR0mNWbSyN6FF6lREt
cm7EuQ21h/R8V6u8RwGO5lUEdwCF/Y7UWG+gNMfdN4nIA5+N0vyLwj9r6bQyJw369IY/tNFWXnCz
bP9bOJvI8MtHDNxSjRHkUreEd+ZRSazCVMkPmjpNJ/8F4RFIFGMqd1up5d+RNVr16DLaH4whb0H7
Bk8mPkvgyBRyxMBbL1W0xza6ZzeACOy0lubcKyboY+Gip49cQFF9ogrwlEh9YS+5uBN22JfMv+6M
a+MPBxj97q+ZbWPTJRYdhOMISTREKAhX74YHJuIPGJPPvag3OU68nFKfavAc05mbjvNlPiZ/0W2I
pBGa7X5gUW6J0RbltNrB7dFu4jb2eQ1Vq4KRJ3tfK5mT9iWWtItLODI5x96VBllUWf3qkRFzz2GM
SZRbKQBgIE4AKvUjp7p5CoUTgkfv8sFQq1FxlgJco+ZbSPVDpPdxP1qcU8VTX7OBWE4i5W7iBk/u
jtV0xzfidEetUV4SgcqYrIaUwXjI2TH6eVZm/bvddEb92ZsId1N2iLjPkirSPNjut5AwIZvPnhZU
RTgBaRfDOfu1u6dZUbTxhknRmwel6V2/GVNnUxFB3rO0mpVFYry8Rx4wG02OAEs/Eewjqt0VX6os
C/ZGQLD+HPhnDNZGMCpnkm0aWx0Nf+dY216TKl80Ch9dV13E0/zqQXP35pwJRnev8raM4M6I7h4C
sh2mw1EV0tfHpdbGOxutrhwQ37vi+R7ZmcmkUVBIuHfRty67lyxYaYbriSskL3dyhoyPUV3lTzlc
1AZ0iANa7PS0mqOUEUOFv+vDzUg9PyTzYClo1gQKSxvT1RGx2J6CngKwWQuDmKRi4fbmFqf/x8AG
jDWCG4Lt4EVrmSBejJ5Y0tHiF2/k1tbK888NcpSWm6kellxLhRVG76+lx/Rkfd5gYt02HlEBYqiO
8qAvs1jidbpacs7UM5xox58GYORAPM+iFocduIC/dN7O9bu6bjvcTGKskDV74zRhSAQeolMbP3sf
wFe3qbXn9NmGhDjtPRFox9WdzePhFHRasQyqXQclBnAB0r4XCjz5Kmm7PygUkVlQMAYEdhcVFogq
E3i3EgX6s8Mrpv8syeMxAddjJhIs10up+/5C3oIVrUb8Q528bu1B7Epg7MgQyfDdNbQA7tKnIeR+
qyBVofLB0FLs5+1EbofZwRF92GiJ+EccaX0sAiA6XgL5yjvnCzASnzoMQuvNXjQ2PA2LcbHqanW+
RmxHvsnOqsqxohAuCo9maKoFpAkSb2okicU5WnUyTR/Vy5tjKk1GBADJuEwG9hSh7r4gLV2bfrUh
dfbnUt+bD4lt+3RTLEvjDIfeKZp1qcu1h1F+cISz09q10b2Fpkl8CEf1+V6b9s5gSN61crK93V8J
dVwXobXwxJltL7HvRso+n+Gqq8UzJggS7QEDu001Ta8mdzuZCDgNPxtzSossK3s7i9+oPXcUIG/D
w2rZEIIGClmG0ZpIUUubnOzBkT8FY91OmudllFo42Bt9SxqvBgsxFg/PLXZP2AusFuUKaj1OtQ+b
ei5PwesFO7KODcW6QARr2i0M+CMag/3f5nCbOqG+QOxaLtru+oFOrddN6bo8R021j+pmhlTToY0q
Hwe9Xyv6zjWocsPzPnXdi43VvZUymOb1WiG08tdDs7TXXuwPcNYYr4wlowmN4IN61bn98tQrhrNs
ELHYrI7bm18nolnJ1DvX8ymITUGRboNEVXRGvSwNL11V1OzIsC+NFelFWOSgCuyDVxh/yia0pFV0
qrFF/o8kqIoIcNDdjrnF8VK9FzCJOEcMWeoMQt9UiqeIhLcNjg6oaP6F6v+fIkxqgt/d+SvbAxW1
VZcZIjShWdRebmRif5n5yZ4qfOqIBa78BhfeiH3BGbJcNe57kZqPlAwqZ65HiFH6gZMo8xC099ez
ujvdC34nurOShP4YcfTXLqTElpviuPNQmd7sPGomOLOqdsKldcrNQhYi7GI7HClYGB3aeuYTaRqx
+uf5juV3EH2vukBOdIIEcfXWlwws/0Qk5WTx/Xj7pDzo5Y4mZAUGoDR959ohAdbFqHgPJaENEIQg
xMx30Q0XZ9cFDtuJ42os8z1LltknARFTvTZ1ynS2XJ1o98mZQ5OIGLR1cFFqnOPuocL02fW7qxNj
NCXHUcd+dg30U/UbyduWAY9LyBJ6bQJrvjjJRF5rEn+qYncEOcq/aVvVIradQ8Ypq6RKIi88mcJO
JB5LmHWlL71cpHg1wjbyKYr+CYJGq8hIa2Ag8pzUpMTXxefmH7QZXc5ktcRkqD15F0dj5gehOBSX
hfX6MQoLJoA4Utf3/tB7yhA+hhsyCYk4y9fiwD0XjzesqRlTUMcklMxfY9z59dLBc0hPoqs5/gKm
A8hQug0G1Vhm29ivlGDFZ8n+r6UU8FVllfEd4Lgkjb8skuDvPxtPuVa0N9mmQfPFwGRkaJ1uGtaK
91yg7e7vf7uRv/Xbj0wybVDO5P0G8zrYVPk6fTOd4nISpRD46BwT0avqd4IBVmKj5I3hmxdBuki4
BcbIhqFjTWTQDaz97EfcurO2aikCboId6W/q/DgpBj9Kv8hqzchSM+4uFSP/qkZxT7MX3SmE5QCp
stR0o4R/B9a9+VTBmp5Zw+HLCL14yxkk3BQE6+2iQ3YXXezoseafdpTWSxBIZCGQN/87auHbPwvR
moqVe6K/tl/TUy9HboNCtNW5yNu7QbY0RJxOneMjkTWafjco9/1ONQ4m1P8q5IhrAVfYXm4gRewU
NP8lmtlbtokNrztZ0AeuR00spUjdCUP/ATjwrq7advJ11Fx1ud8hkAbbyDImVqfwz+9cnvmvj5YY
VcncrUPa7selcxynBx9l8jeuLVwrwtZPlqBwi3suxDdPYyq9GRC7ho1LsnBCAxGTqNAb1u0kA8mk
Nx9Z0Uh/WOmmnTk8EJMVBS3TRKDCcgLLScdC5C+w/VAr68q6RLcJsvSg9FoMe6heMj08vJSXcRFD
e/gGhuAyVl6Z02ke7BF2toxe+/nMn8obgK6Sotg2qchXEZ2V3MzdN2x0rZeeDOIN9w9nHpJ0GqZb
Q6JvIoZnFNOORc7YJamyu2VzduhQawsTyYVZBHJHsxtPcSFbhLhhiXhsCcOMsas9qoCNYhLKhXX7
sr3/RH99wY8YQZ4Pj9EFQA3A32T3Gs7lrV3s4wf9MTmXNvhcJMA/hvrOO4PMNYo096ovzuq1Dc6E
kN65jdr6QKw+4i8XLOt9OBJ/7LDHKL7JwPiyCc87Pj3ke+9fJ1DC8qcnV1RjrkTXHBjckJgND/vz
qDdjSUoAjYENUtnLd4N/pyTBHyf35gpy8hcezKe2C3/LjtwdqyEQgm1RGo7/dnaeTFKuf5tMEgmt
CFcFGeruNRBST1YFlc0M/uKrLt8gtt0goP2PkC/3Br/eb2SpMvrUb9vw2a+mZv685IPWEZVGDz8d
tg9razocoY965WxyCJ0EWK2xgLd484pzL8zy0khObUcHtueMaelfJuXa6IdAi5CtWjS3/viy1xpr
aSlQRUdYjOKCPUsTud8w+UbPLE5ASyJ4fxuJWa8xU9q7WaXjaLooLsLFN1a+9mkjFDHCENU60Hxn
/f6HckLu2dpexjcvmliP6qNaC8XIkAzJOlxeLY7e2F0pVvQnuBoo3DCWwsoDDjLgCZrF0KNSHvDa
4v9MModILi5lETO9suIRVyEGXH69mbHv7mmbH3ufV0i4fJInZQ72gBjD8VIltRrlFGlMtTQya316
nUBgkp9Ia2ZB7BDm/sIjwWMEpRkUhl7Jgjxqid3lL1TGjUsJkKmoU32VunyX3QXWsUlX0s9vtY/B
OTcRMKKef0LXzhi3kkJpaJejD3xm3Q7+x1ggqd4zTIzr437vmLB5nDqjAe5CTHvMWyyTU029R9BI
zIE0dAYakpSL6uZUwVhHvR5Hc01E2qxxB5jaVsk479X5iEwyUltFxfD4FWLxAdMSc1swryatZizR
Hj0E94of4aQt2F91UYZC0iD1+n2IxJTXsekZ5grkdfNmby/gS4VfIJvaUt76IgDKRTjt0LLCco1M
YUxRkqBy+Kcy0roICYqw2nbv4/zyLt1yT7/IoR6JoZ/HnwFZl/qMlx4ZecmY/jk12c9KknOkg6EF
iMlnWI/C1zdSoKgjZPRQhvjTNj7AEE7VbKqMJbSilFY34RZANE50RqEJZDSK/ibSBfpCbfO81WIj
kD5422t4W8TSm9198ZyaWEe72R0xrCvBtzIfG3wPTI+zE1vX1bCr9R1TgleP3NGPqX9gL972kaUh
IKID34df+HSW5ukrOV4EqZB5EIDP13UPp0Pe7LzgrQ9s0i1LAJGtxxJ7ZOv/cKbbkpxUs4ENS4ft
9gXsSwUznSStah+NwDkHmyGreZNBMNESjPwIInVVEoORgcBYT2N3sQ2mXu6rRLeE0wqAN3r1ptHU
uGqfAwGvbSfbccanVGAJ5b+awSGAxZ43AI8blrqPAg77zQzvzCGiuuOIPdptTYyNqbrtQj8w/gBj
Uv1XPcPSE2ut27rDMI5F/wabPYFC9YFn/Ht3atYjDcIteGKsdBmkmNRALIDjaYfbe/iQRvAGmsFe
8EbiEWNYYmYx7FKYXaxL+aldTrajy8Ql1rrGfmD0W/ejlyhYdck2yOJgJC7hV3xQ83HLVXY6n0bx
Pt9QUc4F40E91SP0rUnIiYsygRStKNHoRKsehc6XBfAiUNvo0l21wOW5EKmxGYNmlT7iReWMRnGo
h6bmIRfAw5faNUYxMCIi0Vac+774E/9YDYxJzj5hMMhsb+RDtlULi4DUciYr3GDzuAxWeOqcW/2G
mc1mz0wVwjw5/zyGDTy9NzS1UrlEzJ+xdJWvy8M9KWg6mXgAV+P2aopY+iHOheZ1kkqpMjauG/Jz
Ew97JOS8MPA7nRghm6+vkEWEkmbivG8+rw5lVaoTxirHM/lWy2xVLIOs5UwFShoXdQ0mpIFwwePJ
tbMNa7T/cBr8IBLP5zuhWPiygycAax3rCnDfQyBupcSMOHANGkJCXkvlo1mPWX7BGei6W/VCfj+Y
6Xa665DYp+r1ixwrApZtyxXFB+WyM2uoFjzakbQ56UeDi9l8DHaX/Xd7Kg8NAI0K+SrrHdStCOmJ
oZVIk6h0U4lo9R60HhPNoMCokxbed8n5H5ZJnROJpGvUOUaTAUjADG1XrJjbg2LuGojrqaiSbljk
LjBATGVowg464w6zrjqBpfgf0fDACMRRFI2JLWa+Nulc0LcI88/4qgpH4culYxxw5IWQGT6U/5ah
VUTiOhoA+MOkUkuk6c2F/Ln10yaFIFQj7oWC3vGlrLfeeE244S6hlo4XTaZptUZGHoprIxtstjNP
c7U5aALOIsOcPDp4+7fFI3/kyn3439w0/3zcbSo0nDb8xums1uKhCgfh6numskdFFAbW6yascWgk
FYUPqyRFyJDC2sg8gZiImBOD5m0/qzvahX6dRj9XbRhUuHaJieBfdwagSJjG2I99kR5pQPfewZL9
xFTTuO6UlIumEmOlLR7GiBoWDZo//GxgpliLFjgU8u5e8DkwaUPjzVsjYzbGI0EYEofw3hc1fuy3
37oY3ikjWpRRWSPjjWT7q7321W3IqTnHtM+TAh0ZUlA3aBCeihi032BO4YbzxgtKfX2fxQUA9J5A
gRxDO/rUo7l25BsL3wRFoRH5CK9FQP+dk4DxH5rpLduCf0WFvjjtUElKgZuxBrCIA9g2XJF5zP17
eSnNqpFZ2chFfdL6YwtYRyKJO62VRv8CDUv/aqqKoy7WDBn21knPd3jIS14KNIffffc+kDQHekaO
y4/KXqqEGgzYLAUeb2wxcPnFm8+/0wz7C24wmXNOYxArqpJ19+iaMcNihDX4I+h2SNmzS3umuzh2
2hWzjw2/E6Pwge9MIz1aGwjXxh4XTLuoNOEtbDyNMORQ0j/7x9/936QQjN4lMUy1No203o+4ZvpS
3bqrAUPbia4+F9lUQiRBjg6cpYOHrARdFHXgw7/oUh47S/qPacjo1s10r0llhYXaObF1fL8t7+Kq
S0HXUj+6Cu0AU58deaX/PhSEIYYegNV2vJ79r+JgVJQ93NJfiqat/uFjKjRaPIQIWUqpq+4l7UxJ
V+a7/WO+D3EYUFq1sEHleXsi0G0WKlb6rLM/oXjQskfnxcdEb1im4xzMbi2LDEL085L5al2BvDXz
wqoMKBT5LbSHNsGLlFpxNVcXtSdw/7NBmMeg2qka1TDxiP9sA/579Z8sqnUKGsWRqCUmJjpuVgzH
7KS3F4u/QKfjRCwokTnVfAH3o8WE1eJfxVhUBxyj490XM0VqoxgC8vXKwwhx9Yq2sjcxcA3XUNQJ
pdAYWaYcCN3ZpNSBWEoLy4zvMsuvRErgt5WCw0/9t9Nns43/DfjcLchHlmg47cd+ljT7s49t4/Ub
4Uv9LVxDwYkxPMJv20xt4JHJt0tUWEevpp7eg3FAQPkhS3+UUqtPdY5edFcHYVFBkfM5nAVNtfpC
ADDpSJaBsFfP5c76h8U1xJZkNMzOHsu7Z7mDChhQsc99pVymGeKvxwdx1+uFzRPBViv+2lRa5KmC
fXsNaOI0Ecqgg7j3qvcOOLPHMWVu4Wzki2af7WbsKEu2r3dmfW544ezK+GcTJsAG/Poth76+imBA
R74IdmaCcRqNyBD6YVcmsGsbQgpUKQWaM6jdcr64nGCASfuB1HQcXle3GEPivFTYXYXlq9Kf1MOt
vsw8n365EzYQW+KG18Ty4w5FY4Nfr6VZHAO4z2L+KhEnFsRLxWs/bEzig902PpgZVwbWC1F/eYdP
Wxu1IObX1cUOirXFPXmcvw/osTgY+GF2njhVBILB07fOPrZtQ78MGDe7AKX1jfiuYVHkZ9HIN0I3
itM1psIeRBKkkh4wpgv+VWx7pDkOfVz2hYlYmKhCOiiDT7++NdA9mVv6LSeKZj/8aHma6d371w7r
nx2VxPcM5sHHVDnB47j2ECSiD+4gB7AOXSqhqQkWh4dqBVrqKgy+iqEJqHFXz/YQS4lt89G7+5cx
09JJuC6XToQpYKfYse8RZhDuCpoBMnMTMwN0tJzGczD9L8xT6yAA+Ng8tTZfXCvUlqMoia+Ta0Uf
76rNlgXxLw2Sf8KSZbPH+FeQdSp7hciDh2dV9Ph4flEQmE80Sn2RSZRRScCPar2BEDRB83tLXy60
hxg2i55sEl8vzdjCAusNP+rHGA2tlXTaamRJq833b1lIrvdPdaWh4ecW20HbEHQgz+v7uuYv2lFA
9jBYo6E6WAUFmizh1+CyuRaIBNY0ekS0QCv3XfL9orVJFMxiht1wgA5RZqISVBhiFGxOCM0TU7Yp
zWnWAZyl+MqaOdk4WtNz78Riswbji/N8A+sMKZ+RFf0Wn4pqFKgoxXvv9TT++e7YwWEMSP4JOgjA
i8MKX2F8GyIdTjy/v1w4rViYY/V1LCO00OKpp51MrdelJq+pKpG/8QF75URlRfYPACgXmJRiLPeD
ThSR3r/qsNDghG3iOhGpG/ud93VTu4vyMcLer0Zaq4OoRpAwvKh/dIOTE54U3UEHZ3eoYTlVF5IS
l2rM+Ibwhqzo12CHUZLxMr7bsq2t6EwnM6dEpedmr4V3zFhmb1k2XO0cUN0UESdCN4LdI09ELVvH
Z9wr0YEDzZcV0rebYHqpgiqJRxsNlgSO/KVgtSzJXyQ0mKr+UUzk7EISDPjVkC1B0XJ6GGUO6wyj
SyYowXCJsbVWZCjsUnZM1rvpE1/GzH81Qj74sLzvW3Afs3E3Csaq05sf3qlepJIK83WUSAXyNdUl
CB5UkONsT9j/iMdx2ON8YfVWq+cIDI6O0NzYpkCNdXGKCBN3gXgrsK5GfMBC2KWYHCM41YSdKit6
6cxQuv4lHmihoMCKRM88qpRHfCJ4OClQagVYPXg3YzWcTNktkuXpGCnbWDa4l+qcZS9ttIsdm6VA
KEBWPYeuxqNHKw7uMg1VNYokf5sWsywClFYt1Xjbn4RsH1btSg1s/00dJiZii7F54KCEOoR9xWqv
DyFOvelk51OvHmMcfabM9C1EoFj4DGBmO84eiMFIvV10FpCojdZ70XRfN8YQ8w+8xFkgAlfjF2a6
DEmtPIqyWP8pI3TxbVYFE0PANlus6p56UM6vd7IGSXGPmt5a/W+d4dbrXPQa2t85nUES+uqKSBR7
aRiLNNJ1BMMP0TiykyoE9kKr4NOrTgN03A73iD4G4e+yxWHOzlVHpA73mmr2WOpcdWkdwhWq0QzH
afL8K5oCiJUpjDFvNQe8fzeaaiKb368iXVttGhh2BaS9L02l2q3HKYyD2ZiZCyJENR9BMv6m0PVe
5gUdpgVn/gbMqxZymE55vJjXVMw+PToiNOOl8NgQ4bxrOJ56bangL8Yfasjy1o0PIwXRReeqzGp3
Nk96of0r+hj002iGlBeGvwRPd385WjZyxQIc5zVmj2YIEs9WDtvkKSruouQnfesSJYWBPuTiPNie
u4BFC7oOhSesHhWNdmznyoizFBK2y0IIbjoemCoPJbopLqe1LbG23JcfvZIvL+DQHhEMfAkdqzDi
3rGq1QjHKjsGDuxNJAgHxWGdpaGIWXyZ4g6NgS4GnJgaTTa1lC1/sKwXdJyOkZzXqUabVjoP+fvz
y9ZOCvfqz3P+DL6U37u7XrEabeqM1/dAQTI9W7lhs75zzEnTxRFA0xiZk9vI1hcSYAWl4DdiWypQ
PMlY+GS4LSOOCsI23r1MpZKupxGn4WawE72f2BHxhFnuwnetP2FeCu3sJYd0hN/3o2zSP5AuoMUO
Ok6WMGn5THSCLZd6rLcuvdBwFQW0/lLRD+uVWdqHm3ny/5Ls+94dciHThgyILL0+55k88ruQY5ek
b8kdFwaXBIzhz0xrMvcTM0UqXV/XOheYkwc2kelZ4DRCiwwYdlYsjzXeEBZ/LZoTJg9961o6H3TX
mI9hrE2aqAablG1aPxYSwR8VzORr2BMUx3i6//FYmZz32jinfYo3cmHa99g667oO2+HQoGqg6hlh
nsF1I5yI/j/vB0HXuwCJXixjItHqt2rz3BSESAyrTOSUDKef1fvBrhTS6AAnzqcYM41pL/kDcr8O
MpkhAyMVCq/jVjmo9ly+Pa9kVfMWTj6hVacNhsALNkwb15e3rJbltvgr6oehyLRbZHy2NQec/0s9
ImVz27p/HjUNpsynTP0OuHt5W72EdFjL9mcWXhHtCkLYgepoQIXzR26Hkw7V8pJn3pqiIzRyGAPk
9LgFhFeZBNkmP6pM2vMdiEblFzh+yBR58bjvomdI/sIev4ua6o6mVOBM48RocTxDWUHuoQUTwIoM
FE+RTViXFTe+q1QRR87MJRQPTJQe7FsTPNEGsouqCdfemTfy1OJ+s3xyyqjQr3vjrvcHzc4nisP4
rjFtVWhXHZ4X8Omq4+IWwYaEKUk+gcxJs4zYTSzI0c8Ulu+nEgvX/BR1z645nol5GhPMX0OH2Lte
oU6FlgwVptYtR0YwaQ1SHQjmHvqbZqF0GZC7axKQZhMAUzk64+sBV16LS7TNpGJ0EOv8CF0asEKK
gu7ROxeYa8TvODqb34CuqmP93PHHD9yaRqsrhjk+d5UQ/TyVUVdi7jYac6alnORww6OHSbtIajXN
WIHPtZ7hxHGTdb1gT21CwAcQBxfS38WOJ9pUxn9QkmL1nc6rRA5YOAGkVCLDdfp/PNGgBLSlFTkj
zr28t5JNK6eQujTuE20POXmPQxq15acwh6xeSxu/Q3xMEGWg1ifOsbjpLZcFlmhdrpecILsZAVQP
juPeRtXOp1yKKUILNZACS84VfL2ormvdhAplqHbM3tZPKUQPJTdLVBqINeMJzsc6r7YC1GY0Pf8t
hZUlGeTM4K9BZH0ln9ekb/p8xlLHE7kg4YwqHuwII12nPJPldzQcxodsyPbgpjOgawSYUVobDrwT
qDdyomKRC7vI8g1yhfm1LEzx5ldobRKydhb5TPBLqinPOHYwUrFYMju30mNg889GkBAQ5d5sNJ67
OpEkUcADbZdFd1LApw7AvWt04k9+ZvGvjgrZXpSPl/EtwteADkYgO+0bMkx+OQ414W0oh24Bzp5E
w6N6D27N8godCsp4sdgkWWuUzKwzU1LzUAgR1O0Yfxyqxwn/HHD3XHOGSSjvf0P2Mv6s2pXQ5/sS
kb4zsDxed9VeHLROwCxRPCBhKJdD03y6RtTF90brGRuYZ7vdY2eTimgN0BypNys2+GQKXkMaR2kt
bUeRYhjXxIgKNmTr0TiXEgIyzDqjhUXGblmYsYHSotuwQmRXfQhtfXrPbjLpz9jC181n6apfyFBc
kb3tXmLSw+IQETt8oecI9Xgi3dtyptckbVDEXYV/5JAst8osBcydSUF06c+YvHT+LbY6TiknWUx0
p9L43W1h0bCWEfFjNXA1lP3qhuthlvMdmRJmt8N8JbFnhqNGCIZ8N9G1+5fxC9tFN+8fnl8uJTdO
1ygMHb+6ThxMrkw3X6fjttef+fR8rgO2bnK4XXpQF9ocmmESh/OciO0tVCOUv0gbFRxx5ESugEFp
/y3T+pWU/P6hlzYX4WTdWRVg27QvOsw5O64mzv2RyiLEJERD9pN1M970SkRAflJE7NVTxq+JSEkV
H1hMgZosCyu0M7ekxAa5jCQE3mYMsSWNx20XjJ3cKqAWH7kzlAVMkK20yPTBrF1jJs1nPQVn0nIS
dFdrJj6Qm+S8lELXWv8AsP6+Jhfmi1DTqqmdFXrA6UdIx8m//cmR/haIhOw3OjVywNzynMChOHpW
77gn+DMZzSaAAt03E/UzLnrf/sVcWFZg0PN7HDaVWIki2GN/0R5WzV6vKHfL176mwn7ES9oH2Kbd
B0NGe8OBe1kJdIihu5Xcxqk934sfMgJaEbtufUevxGLJmraFE/nbsNQ8fiN1ujA4OsoXVcF7gJqs
PniLjjfIClAg2CrKKtSGNGpICsbEzFGLUF2Zs5QQpP+pIsngKqZTEIgs928rddkKW/O41e2JqmqW
TZXQyl+TcMXUHrDo91dNbxMMyZcjFj/0B3j+e1FGbS9pYy/FPXhI//OCiKB0x/7kI+ZTeDcZnjKr
xvLgHQLZ4U0PDG1hokt5ziPP7oLSdGuXzOV63ZxobZWdRbuhjmiiPRPohIIXDd/1rFGWgbLhJTM0
tYvcsqpKWxy24BAaY7luqof8jLlb4i9Ec1SJFCgK5oRPVVuXiKWaE0L8MS/7PfpFOrTqv/qpUreN
NLryaAFLXiwFYKJAx3trz2+Vr7XQxDlGPzD//4rsq7EwHWSLjV0EXZTh2tc6ZHjUyq4YA5OGSmSb
ilfF1+yVWILQwrJJL5LilDCPpFMTn2EJunuCIY/xCL0spMC5CgS5yzVYJhiNOKe+78e+dqi+Byqv
Rek8Ix9AXJEEgXxYZTRBoS40FW9U7wSjuxW9RQ65IZjpbBL7Hzt6PdDX7J5YEHN86s3gj1eKPUtD
DICca9hXE853o8slgAjLIz3tFu7d7KuievI8tuMZBE93W44hvdIoBZcnIfFv2ql9fHhz7PaBFF9X
5EWh9Jy/832VUimCczPP7xXZDIjnFEHeJaeMfijIpn9YwR/G3iUBwfRkfiGbsEawzgABfe3i3L1r
aIhn1SsC2nnH7QL1SaIDcn9HPtxj+JDlPQF3GQ3odyV48H1unvqi1Ze5nph6aJcnA5KQ6ojy+dYb
vcKIQQXR+UHIwcgiQlXwmWki/hn08arTcLJCld5DAASXYxObP2SGs1VWsfo7xWy17yG6Iqus0UHf
RgTM/XwCEx4hkA+4shyDe6o0Hj3y7UCl2bVDlycskCHGxNIbwmz/3kdfMQxf2Ll60CPaRRoH9FsU
Rjdnr5XwSohQTLGfAf/AQ+Fv2cmEhUTp8JPMrtDoqU2hc5z/HrGHap0XtOrGtjgrin8L9q/ggoPm
gCJo++0FBPSJ/Y4qG/Oqilq7xSElY48hHFi/Q6iZkV/uicSJY0QSLZpcIF7CYscmwtFPIkDDQPpn
+4H4dLGwWN/BwvCppZPxD2xWey37QphkH3qA9SvZqeCv54z9lMzH7ArDCfDGpbJcT2SVfP46FaGc
bt5FCWPMRvJMh1r0ezNfSXg9ED+GxMqkJ8feVZKxK/9dlIKc34tBI19YQV9q3HR4Lez508Q9e0UC
yTzxwnjUEiw65FtVZ65fksDI//qytDRw4hmlEFupF7I4gsomKAieaM4KGdQXt4m6fpt5sVzKfxeJ
PrZN4WD4Xuar5UcujqZzUdmnn6yHncvU7din8zFyYnnKrNimVy3RXwSJxgEVlGIltx46dc8FGOEl
SAmtUp0+iV6MHJpxaFgHgvEGv1eoVTR1EWw2nVD07bZPLdD+kNFE5tC8iEqJGe3VSrJrj21emd6r
sXYLxspP1M0io5d0K5wgxETB1NphC0Lc6AbwXsr5vjkbPs1YuRw9AEeVlqwZLF0g8BK8xmibOY7S
TfcGFpMSCU+RvKglNySIX3r2AFmxOOsguPn5RYsL2Nr/52ITiZeoJH5JVakgZIWcJsxtnliRCCZx
1Yejug+1DeWkVG9jE368IW+M6+In8KJetQhpdeh6vbdoGAIgQJUo3n4jvA6mhByAhds8H0QTkIWm
NRqYIVlIS77M8jcQ0s51WM32jm+o/9eHZhG2tHebZf/GJa98WYKhzFk8dgjnZufY6ClMqbZ8LK2S
xelN4cpflSmTH8JF0W8hEmsghQlTZL91Hzx9cfNJDxNcU4a+D0WeBefJxlmuGWr+CIxF8V4PTpf3
PuVr0+7/XrPUKpxkDB+ECdjmOVHhim2C7Gwge3Az8Z1HqaNc7SMmje2pxasmMwXzn+MV3jLm9uwh
fmlVO8WJy5VQQGJaclEFaDcWag3crkQQ1EWBTtuRqL6ReBjaGRBxjT5fTjr+5AHwyagl5TS15JU5
zz2mz7S6Bp0N9sjlrFID6ZKV3mVqrhH1chnoFIBp9IinnRisymHRE/713oPx1w9rQmdpAViYUiQd
Wsjv1kExKjtGwjB9T5zLmhgZl0oytBTBXCjXTfZi9nBI9G9ZuHVWCAUuCB0Xsau/dX7rHlHsQiup
qVXCMd+2/4igXopZyGPSEFlG3X39ds+sXPeAx+vJTAC8cvp/TFRhw1kc5kn/aIwsgeWnDUGoMTar
qY5eiFUJInocLxV5q9d/oEFMFc42O8CjBxPKZxR3E3icCXNx21f6e4TOXGfp4r8qWA27iPrwfTaO
yVR9AOGvD+ZKoCc2lyolPw+Xj4bnQ0KB/mlRE7FZucvsZZJ2JMCkB1I8eaJlmQNuznpJo6zD2sgu
+MzypBLpJJscKYkx7RgLGclQLPJYwWdtCOlD3KZXwPVbtWMVnvZto8Iyz9IhX5+R+Mg97AZza2dt
b7oT/mOoQcs4mnFEViUdr93tX1VvNyHOvhkHujxAfaidre7rWC3IVMEj5f6fTsWa5b7fUYyQ11hB
KpRW9VmhA8JvFcuFtTmPMtmDMST91k5bTbbcrAN9KDwLj2cXcK7ia4K/LoSthOn14wtUB61v/4TZ
oMgSuPOC67tFjuv2i3mWt5/V3RFAYTdL/6f3lMB6HWRM2dexj1P3QSxq3DDvHtwmig4QIszspXGb
y1+CmEmSGTSgbtmhAumel/1mOm/HJjas97SBNwAbENusuAdqF1T9qdCDTKiiPeqU//GEHIZot1Lm
XvokwH9CwkbxufTdauxgFWGAZ6LTOJItptnVWPh47JoWF7Y39xjTmu0/YlxYetjoX5miSt7KmJcc
9YjnsqJS0iLyS3LgCYSXAPKjn54BZdyMvMvy55MM3flL/MjGqBaHUxeMny1sh+F+WrEpHqvBmDdy
tcuZnY/d3+P+rxsqjU1Xh9MlMh4SIIlselWSiCwpvwglpMNg2snI8DlzozrXF38bynOyzvct94bt
x2P5lLEGbq5NBBvvXYwbYP0R2pQ1z93mzxLcsz9lu+Gf4/wVNB1N+xdLaCgyyfc2AimAdQnJTWPR
mr7n7S5YejEjUCEbw3KzP1Gfpc1T0cktXMY++3jC/yKc6TjM1RhHVZzdoLae9EZrAFvk4MRXIvX+
zBeEWFgfVl8bIuLUjC89128i7mmexZAKwuCBlL1uYS5rjHHWxzyPkxeWS7nbVp3pXDyfFJd53rP/
WUdxy8tOpghRudaNh3/6VXCczEiKfOe4geGH5fe50xi/accAGnRSBsUJpHUuM89cVkgYSzFnmgPw
FJumjwbgnE5U2FhyLNvfdaUGhfdPLGFc4Kso+9vdq19TwBDCXMFMPJO8xGPdW3uvIpXpzwdDlne8
yGiyOrhvIJZBDVFp7UxgIbQFyZvNJPKDMsarPSXpJ3o009uA2C1qPWLY25+KlIyqOlEYClk6HQWe
8bqMhi/q6VIryk6zU81va7ILTdEmBDqlS2NugdpAjjVe5JFpGfTsRAjJA/IBu9F/V/nRICPcdFPG
07hqNb7uGMuME/5ToKLJu6rFUalhL998OSeUaQFejnYgwFJspTQVaP3xYEyomjX6aFDAPPiJUaoA
ke8vpirkFQg83VqWDYK+zW6lO9hDnhYYDvOkkwAgbEFPDoV+b0Ub3l6d0NV5yGMsEmmXUVdWyrd6
iBehs2mshlFbYcyHXOoVUehGdCfQWEKrHE0Vy06uY/xvR5x7+O3+WC8xzlNWMevx4z2HnbE1tU58
Y208kYU7MHMqQC6Xt7SUYwUxU/vBTg8I+PSDJIQqTJ2NemiTwl5bZqvF8cWIltDARu+88/49Fsxe
UnPw8DuTlPSwhe3CSkRDkUzNINzVcPltUyEZbJgi6yUwBIbNS4TJ0LIAALHc0SFsFIPOFCvOvUzk
x4J18vtNV7V53vg4Ou7FjXNa2swj3gQ91MpUp8g6vwEHv2QcK1o4/CaJEMGg3FqX1W46u4gWJBW/
hsEpiC0rbOOAkKBYHFl2RVJbKnju0jjhLgRXduqho/tziJzhfb86jM+lZsZWkHk7PUHWrMJ1lwPP
LKTaXWZ3TVET0jvMoh7md/p7FlQIZmxRvYxVdHUIxPEj/XQ1RyBiW6Z72Aqd3nj4DhhCrpzEL3Cl
dvqCmYZjTAvuLO7UUddlHS94uVnAvVO8uH9is/2vTZOpZ+YWPIHGpyeghNufXWSMj8mv8xc0w4Er
m0KMEpzmNz6CqJY5HKCx2JDrIhFqBdbkF7DzmZAg7QXTaGlNZJarPV8zEc0iraK7JZICPshbAbm7
mx9xHhGfLhKV2kqgfTi2alKRje/Zhes4xNG2TcvKdq0d4vmu+EK0pELPdftzXjgkNDdNhNJiA8wv
4sa2jcq08/S+nP+GewJMub+xs0ZX8q+KOhuqPvdWTwONd/ru5LE9TVjgZmcEFJz9QwvEdXYe241X
lBDnulZ/1lSh4SHn3YiRdMwjIrlcyqZgzHBSBcOZgTy5Zqt+sGEkPYYQZKflwqvoiBs2lGWDwe+b
NS6tMms127YUxar+bXE9NpxwGyjbmS3t2VNJ1+UCIbjhsbewTTn77d/MCdKOm25XjYvzp0sJP78K
T41dGorzntXOxDpppHzuGqYRZ0lf+sMA4UI8qjB04gzuRaAQpqMN7NJJYkymZjerVQuDWMWfcYY0
TFPRsHuee4nF2R8f+sgI+J/8iBqSK0ApnudBKJ5WQtI6C8toyBUvKhlSOTWAyx9mSMx0u/Q03u24
mjTNFXU9qGT8Dpa8gVRtb3XV82K1cFBSVlfrAPhZSUvHP//GUdHWipvxzWEOUdKJ7W9KZJNEOHPk
2twz6fldfAXCSFFLaFR5FUkgG7G2Kde/1lCe8P3v90FEdBu+WJtEcpayszGshMPcVpifiA+CwQrE
OKgLVTQaWenUegwzKukQd+u6IWJVfBMLea1Q5TihfhGKOYD0Yt2GRPc0c8mMuSzDOmWxsywDlLx7
Xb46d7qburVHt40WW+K8lvxYS7vm+sa6QzS7WSt0iPSp7V5E/7UPeVdVyDGuTTZP9cpzdwvAOENS
36IWOgkkk/d7VSZga7o5z/n42pU7sKwL4RXR+WT5YXYLXYEYs88G2jJD57JyWS/W9b0HCXboYQoX
LkajOaZTL+rOAJBLKxr8uNjRPngQURGFYIoWGLdRwLAd1mxMwyJ9GBhQlAZtXncnJcFUXR6YqFe3
Et0HM0RvFwFoc3JZfbFWEGHSvspd0w1L0xYv6Mgf5jlFSrIlo0m59cKEDulJ1SpiDTpByDn7j5rF
WxG7w+jioJ0dSegOjgfQtUGrZGgeGjQeHN8wppp/1oRh5yXYKy+CFIGt1wEAIeq2bZfx2anc4lpF
JjmMtv8Ya28sBmD68I2qOPZNrVZHvQHhMOkxvAqQexqAucTu1SFpnWpK433SahGwlHUVAf4byZpm
EOg4IcH8YsqtF3W9Ix7Uzc1GhM2N0Jq5tOOCpCOrqoTJ+px8oeEJXPUpP+FElBs04Vz6/34PwN1e
L5sUlm4dNJ+EUL4TcADvU/NftrpY1YErTPLJo0tEVDMonH+rf5wXviId9ZFq7xuu20zXod+dStiB
ms6gGUJqhHjLqZpJ3ptTMOteon8qeUEAJwJihIBuyrR9VXYmgHGAJaGrd7Xuv3c93ya/DL4gFhRE
YlWVRwoR+CWoFTn0vHXRtoefgdHK57li1XjbcjyncSVTfLI/KzJc4wKCwIeoWrN8vmlaJcn+rNzc
DR5hIV2LOxYWkKx4FauuozlM/Ab0wQNBSzANhP4RHOgBeQos0jxQPah+6dENNWWZwTHol0vUi+jT
7GOiOkklZfpFf5xTBldBmXmFVFtrg3rQFhsB52N1w6yUKZoAgy72DxkJHw1BQ4lkS1rj2PrBWCBI
oKDUAiq1OQaEqUPEOKHBODLh0is40wwmh+eRvrwg1j1iM4go2YdYYr4Wu0PRXfPNeTE3m9x3YXFq
gfmOhGO48LgoNariWR4VMv65k7+WvZ7HqB2KWaQRfXlTM2WCLbYwC8Yn12SxghTmjDXp34jXTaW3
R3WVSjoEurjJrE8z7jsVZSkgUrNXyNR2bRHNYK8ERg/tmYLzvUmDtgYCdn3hdLhn7ahoYUrJDFn4
PxDbmIwbz853TtrB1SGks5cy+rdOJ+O4T1SFBn49/wNd43QsOA9YLKyoM7aY+4VSaji3yoSCYyVJ
mz1hhnPn3oLYRSuGAgQFR+HqnLrgeNcjKaftWEc4KM599N24wnHK+CbmP+bqEwIugSaz/DTX5f4S
0DH+Ui4Zfg22o9QSCU0b1rpBp7ud9THPbZDltmlpb38hEO+1szHKgYbE2M8IwPZKOcCunJz3QMHC
MKOVeXsdLSg72RqTkyc5+JVSQd6VEjEFduAAlubmcxcJ+1C5TM2Gd30b9UH7nB9TagmPTHB1i0JU
ssiddr8YP6fxiyP5LZi0bSZxapggc/77Ojp1dpTwOZ9lPueptNsuotFZ1GGiJlES6YT1GF6ODohU
FLqa7dir7LQwedqFaVSml1cj3GABrSQ5ei3oy8C5wnLjXVR5tLERQJVwYAALydesB+gVB6CkRTJg
YfdqCEH4rnthEhK4ST0T7FeQXmMilyFjj1Y7fLHE84vgk7vx6DuY6ReCv9tpJU2QhKBcrfzg0A03
DgpFNz9WlrCOFvL2I+SIgMeClezY2mN4MAv80g7z9xhkSXTafZwMQt+IV4FzHVmnxiZd+2YW6BfP
FvPYUVn45hZQzCj13x3Nr3bb7w8LdqmAf16Lfiu3VC7Frc/xFH/HvCLAFfZHCt8yDiRD00GiQ53p
UE3l7SMCW6TJ3qs8s0Q4mp4pVhzzCBm8j8FTBcnUvdeGsLP72dF4tk4F8U+/bGQitCqm8i7CRbZu
/iBqKXj537WcIdEinl8Sm2ZwKHmn5s4FpMooOJCgj7P444WikEV+4tMpBPR63AnTz7Q2WFBItCQj
y1ohRk7cevCFz7xojKXJU7XMn+8c4gs1YV0SBA93WABZkztbhbW5swZuSadEahWWkVtksBeb2Uls
bGDsQVbJeqtjMPCXoKHiNT6Y+DDe+kb+nE8bHmTPygLW5GrYB9qFFPQSkPvWq4+lDFkl4MDdPc3M
tbQx5eKCWBSmFLhbSChfklvBWda4PWQSkYSnSJoDVokzryXdDmTRGLFQ2+oXaDqe5T9bQoEgGjU2
Y3QoijqcAMDcU1tp/EBhAjBr0xGr61LOmqBY1axDskLgGvs5+mjC3owvnQ49GGmHQ0LAqE8h2zMx
qaiz8PoqSNkgYlIfJ0H6h4tKK691UEGrvQkFqWS2G/L/kP8UfAMiVgiYcOb2enOmzJEDzjLkkHH5
f1VsC0p5q3/uAFANiARbqb2iJUXzcl+h6t9d/RptSdz+Z6pgsz9f78XbdOs7xQbeGakI/gucbsLr
QQDAgFmHDfN/1tx1U0EQXNPLFGgbI4GFFPp2ea9uGklLQ7R7gmPUEScKf1i5TXS5dpddf/31USF0
KL/qgh3YKHJKoeFTkZw7eTA1NqY5u+alHoLJNR5zM160O2n9IWGsDzMdCD0Vld4/dBInix9BPE8A
YwzNMWKVqcDRoET/iMSx2X+4yOoHkdtlGdo84qrtOj5qI1N+rTX2ThN3CHrGLR74W0bGFanPSq+g
ONuJ7dXpGbqlpLG4bhnKxPzK/KOK2rTVXCkF1JizbpLYUp6/vWvcs9tvw4TCydluSk9Um4FfiDew
xwQGgFPOaYS/atTCDM2IvDKcphwruYrC6C7/RDgm8zqcH6RATTLZZAPNEe13j9SZvi0YketLJUO8
8LwkWwp7GnZS8eyhgSXYqJ6OLrqshUqydCDFaO87inmoPsDtTZANneMBubqKz1CEXIEOvqazDkPt
9yFKYK4bvFwWEuydM+gk4ZBeyw+wrv0nAfzUP65ZskMb2G5KR7ayMU3C9ZVYPhGBIudMPF+jZ4qM
vnUPyw5D6evOh2aT4Zz6l1TXeosP3perw/L3ISmbjTI7F5WFy2fzuOs9XFPxHE6t8g2QX8i3vG82
EcrI97w1tkr84RT3mlx93SIGhTzh3OygvT1Ljf61RF0yZGCCzfnBuyymxzno9EZR+UAXmlRQkiNK
SoKwjPd5cnC0iaiCjNzKZ0b+96GQD1ePS0/dKA4DuRIvmBONQU/TFAOFC8rDQ75TCxrZ+0gV28HP
YI4ObX9TbjDuyH9279fp/f2jhbLyDPqSnTeMKbN/sdgbOsJtkdaSHFZVVZIaPBG96ccJg5MghaWV
zOu0/BaNzbsHD3DNVT5QyzKjrvmN4HHcTBK62UoQyR9Uvkf3EJD/UTSG44dFgv5S/JWsGpHyWpbs
wqSzKfJhPzUzoXxwfZDuLXsHIZ/XX9/WtlZC8QmDwcmldmDhDOvHGSklR6DPv9reemks9iN8RJ8P
FkZ2WzzqSylIEsxFATHywMunG+FpJR7/MFv90Z8tFlEdaclt9PQna7NefIJIK+wKa1m3RqBacSGQ
fZNnFeD1J8upQGohZkCeQenZ0MRHsf7/5jEWE9ZdSr2Ul2eBgxDSUYAiNEO4ZVZrAXP27BvI4gSf
DL+bM9V5txug6tBaywnV4qDDTZMNn+IjNgjZc5J/NP5AOE+6K5ICJbO4MDA3NQjrtWNEkWcgXQrG
P14KSzAYrchRealOaAa8ZFtxdsyJ6mWHLXBt/tl8l7N3msoVYuMhxrSPhTOPhGNrLhXbMIJ1wH+b
3SihMIq7DbVvsFbEuzLSN0J4cZuOjorag+VlNHsRNQ8B2RwEZ6OGZLj+3KKtXAAZAqZNr3hdImG2
te5Gz6+3Q+obvFFk445LjPG2IS2th8yKveBloyhji8MX8LiHhe1yDaLDl+WgbeymWLIlht9x7dgR
EiawV5msXZc8ZzS+3VDJfS2IycnNhsakQ9qtXDl6KI7ojjtgwo6p8iIvoGf62gAgBJFu6hQfr6gc
+Sf+A08FUuVnFdFIu+7tR0jv3oUIhZJZPZ9TWtiwg+6roS9piXWCdmAnTGgUSGQYChDwI+eQ3qUr
P5taqneJPH5JTG2ASeDUo+O60YTEeaOgjSNLzfvZbgXr5QYTaSseMSPWXVl+5/jq3/voD0OkYiMc
eYN//eyKlqBWWflAbxC30cj2zPjtB/6WV5P0bVdliotLCLNQ5hKylYC0xLaRC6ln5fe6auA71FJe
Qz/UamYd418KNh5yw9R70ChIS49VlZPUi1Ot/Kw55rLgxsqx9UOPAe7RFfnuT8gMOrM6Ce78WKXL
8CbdEjLj1tS49JIhwRpcuS/z6epYymfsvhAotYEnuZhRkAmHfuNKIDB1fOKv07kwm8E0IKEn2jNl
TN+xmPjLwHEcG3Cm87aoijDYk421Sqq0rQgF3wRx3yO+P7FFCYVjUYPqC7wNOOg8+5TD821DvUc3
ix2+AkffDARVf5K1svvWLsi2R0BBTds+WdgXQTXGKo3l4oPP6PGalcTCdNoTve70NfCsBgVvxpSz
/kPv0Klh7jlos+eEAlxTlyjOswSivK1XAR0xsMmnkV5spqz9qslQc66Q4Wz2hRn6K5caFlo/7EKb
M5L2kQmTS/0gLpDQmzkFMI3aMNovZKSIvtEd7LorhVfKdeMrg/zxAftGNf5A2GWSS6oK/wlmTKAr
dkLOjEiMlOitP2El6HI1wtc+SO72LcL1lzEzDyHQcgD6K5paiWwryDtR+DYuSW9N9NLYmiVXnwTu
7Hxotoz3w/OPLnAnNgxhDAhLiyJHruNL35mEJJ+Iu9E4r08mLTx6r6JnZw2UtMXFjaLk0oInfIvL
/08JkbwufBfE5NFRQlB+tItcddWFP72yvCdHv43S6CK8qOIyIITe9y8fTHz4tRbMGzzYo42x0vkY
m6o7aoZgdcMuALPkbnAbb3cqtIHz8DiMaH6tgpdQcHlHkkifGFm+ySYSngLXnzHKmkyBXqATf7lb
kgcyI5UmV3c9QubPJbgFAEpeBNt19rgVpCWkI7B2P/TymQORNcMfCS/9DU4mjM78j5ZOOxvhutGl
ENPnKruT/FjzEYisvFjP5R0oHCfZEqeDuv7ahBqVI3crkjUsDhOIxw6lKEZRSVIHFchUnfMgHTOD
xfjsgjVInMa3pNkcP+NblfZ9eeimkqEE8on+Dc37jBRav3F5veIz4w/pAYxv8QAsMrHLDJb3HSAN
Nh9SFadh5HjkXEl1vlwFz8/o0OLtqgU8lgSIbLZEQRyxBNFYxwYeeoyaSHaq3Tp4lp3+GOm5J82Z
qpkepBf0ceMJLybc3ngSiMBzf1NVrvReK41J01cYdLb4eg+xGzrsNt+DXEvBq+WnaNkHMB5IdUTL
Ayfq0S+OzmjNMQficdPWWfPCvYnUozTyGpOkvGrDNucQssfLH6m725KjufkS/ZvH1JpuGf5huL9g
k09BFdZswJTvJlGNbYFXHH/w8Ac0lNDjaDcVmKrXVhA8vz5KmrxxpKdVM5+Uqn0DT05DQ88ud4+q
lEIWB2i7a8Q0s2VVzVgtPCK1kDUIdHqLIB8njx8WFBz0L1nD5+DKdrmZ/Ssjaq/pR2RwBy2hwqZW
GGeMExYvxLxkDqBBebbH9TGjElN5D/lKVIZPaRXiuVQRB25w0eJ0RBSFpqe733xrMh0NY1r09v7z
cc/Ia0Q30NSRfaRoXqJRHkFUcY3b83IG8pLnrLqYuoDAnu24WXJyq+c2KSzfth4XQbudsbIW+nWz
/pCai7BZ1Xl7KiQGL+WN+2Tauk3zmMHkV90hfxTmvgg1ag5k8BXWL7GT3RK/42d6aqhx/K8+MzGc
B6fs7ym5SAPYKwm+wmJkgk+cveZ3PASQjyhVjJy/q+Ga6kjVy/OTVyKoCN3kjZbRAMx/IybkkHce
qtf3vI4RAyNmVItJk/7hmrb/rkGGCs+Zb3p5kWvCsFC1r8OJ3l3S7Ioa3gWtkwqHTYSx/lZ5f7Bp
EsCqikbCUlZdmTslzC9JOqCnRVlrKIxbyEBSHYphm1n4W4G+JYMeriF31pHUPt8YYJbRVrmNeoOg
JIO8JI6phRZ06Ahf6XUTN8jSPCd2SevQx2Hson/GD2BXWOxTDIdS0vnmLM/J7nhAxCZX3ykfFA1i
WDycxDWA4auVdfPSm4Q41Cnty1K/c8/4cbbDZB9q4UyHs0L2xD6jNYmoAso61TWhXgkP7oHiRcOy
HAD9ILGBTg/UwJN7cqvj6kmioDKDkZLmjnF3hbsp8oBJAtEeZ3nujqMYpu0x1FZAg+mWb0I3b1ov
H8fM7D4qvqsW8SwmTEaluZtSSrnGYCh/Wns5VVslvj/FPRknX7g5TU+Yu0Qo4rqbnaQDLrycvVuY
KesHW/PTwmRI7AVoVocePzi9l3AOE0CYV2OG1U4Ygo+i6/EnJNdai3wXbcGJSAfVmKC5egtVPS9v
u0U6rGU8tAfPX1obJBWN7qwiy7yItbDYGTKrthL4Ci43c/M3OH1oAtkaUJrrorwlevkMFXhaRoUC
a64BXX/eZtrz9jPqqdW5kjBFTfMh6hwMCHWPIFDOASe6yu/oMf3sHqJes+VEZJvOG2dJg/5UbKFy
ZEDuLS15ESdzLN/MyUZmXVUb6CVj1xBLriz4Uj2egAekCLnUkWSAZkamNoLH3Rans8QoBlHGFO1a
xExL6Lb3HKImJxrO7nOOQgH1zMKkhuOCNZIi1cslgvnYT+JJ3KzPHwSHvsOk2pzz5CKo/nAbWTIv
ORy+yYM4Lx7KO7HF1VRgUidMm44AejZDQ8AKmAu0YefcCQ3PIQOtKUj/0MuVXhbCOm5A79poR75v
PtWIQZ7ai+k0LHIreLJ7bi9mFFujMXo3RlEqqP2POsCH/QeFPjViFkAb+R0JtntJUWfoDavXfoRd
jecNIiBDiqpWq+2k839F0DIdVTDSVeDL1M/YlW8P3HtY+EibArVwAj4i9Z/pY6BszoC4+vRfPgia
srx2H/gJhB4hEJiiYyfuue0VzJqDPY28YB1cpmF5B7xoQOiiRzpyRZyBQqKSK3L2vqE85Y9Is414
zljWyGcTIzIAg+iSje8GjBXYKAMqKoz4YTTqPAKOhaVKg64j3I2AZDW+8p2AW4abzZz86ThYS7yj
ElToYXcImHhNyKB0r5ejObdgYMf94dsxNsZawl1KU5zQq2SMYhUQJRujDsl/+NNVVzomQr4oIrGR
CBYtOq3WbYGuOmLqKgaM/4wOo0nCoSoJZUaV2yCipyM4v5oLvfmBU0ifeKCmlDY+UvWD87RWSHOs
28GoHIVpQZhaoh5NAwO6yvi0ahm0wW+oP58Xh8z6USN2YDL272HJzfxITOUxxqykGAwzJk9DeBIC
Cj4K0YWIT/Z+NDYsuQ0s5v3FE2d61CAtWZT2lkTiTsYR+WMkTKrKuGI8UqvRlGZSctAw9R8gGvd5
GKJfIPW4sENZ70fyfTJvGG1WwhnEm8pZLxH9U3VRkdMbQ0X6JUR2vZxLoSkswvYPUKzNmqzbqoK0
qRo1LQXRSyi+xbeSqYb/hZULwNb7pucXEMAMTXld+k6+NhsBoX4/idxuBMh1/C+llnrIT0L6DrhC
X6bV5FTofZhDiSTIa3ZCmSjrAxEEJJxaSztnC1Qy2BpaewNF742qVfHj+gC+U2/Uivamt++/lL9i
sukM+8ozKKnaas7pNo0vgeqDN6Wpz7TqWpqDMjnLorYrpifWl9cPqQXyTwyIKKnHmnEEplT2Wul5
VRz+u2cg4fuZRPLxjYC0K8sGHrCI4R0b6ayhDeJxK03IIcc5tE3Rdk6cwbPZlKpw+SFY4cuYfoAx
nC5GruJiSGiLze+e4xoL7L41O5T1SDl3zipX3eEcRp2xtdVVfrQxfvopMM3J82MVh4nbmgaITkk4
YqrZaJTXNANqXI837LK0AlxDF3jp5BoMPW7ljc+/ctDZ+r6QCRQJfdUZwz1J65goHhsTYAn7TnoH
yIJzG6n9qqh7bgR1pfZvYEie2UdD6yhhPDW7BIjPFy3QWeu+HaJkHVYVmDcDpWgW8otdOfQBKesZ
/AiRaipbusoLm7L5oRBbsMkAi1299d19oCcRlezbVvX/O0KJzdMAr6Z9qJZ+ML3CSy5R5auc2+ci
Mbi26fT6gINvIBwBGCHjZ8h4sIUcPvHtdir9j1JQdNzgmqH5DlkAw6c102CCALVmzoE2yhvcP7U0
Vx3MJVN+ZO245n6cGl2MEvq86UQNRJml/Q1M+Lij6E/8x7ijphdLRY08AVgbe7xd0wI79zPC648z
qJiOImLTba/POi4LHIMyUZ+03BdAhaA247XtrDK5BIAJP5xGQyjfnEUjOcoRUQIQ7AaP7JbF3I1g
F/aT/9ScTd1VsMCsBk+IDbKBnmxQhl3txznSGqn/A4NMSKcbqN5ldc9B8biBK6Ur7PkOZYYv4/TT
c8JzZTzLj/SZHYWFsQsJ4ONIr4z3NeIRUyGAgiHaZV8cOtbcRXsJy6vlp0mV0lQ6GvymhocExjO8
6HlrMXH8B/WPXPGKQJaXcTSkySIC5bU72ac3Q3XtPY+aS8zXDozEm04Kq58X1daDTAzgthX5xsIo
2YvzeaQ7bw64gdZPx4b0vFpA3J4EabQ2Sz5DTxBou0MVCVCpkovfQPTMHVJqaxX4SKJ04IUK7cCp
rXDBLkt+Tv9ZibM1B3FqzlBWTzk7IizUHT6h7CP6QZX16UP2u3LzzY5io2SRqRlKzS9xPkkV3APJ
E81tUYlS93zDn0fqWKT9p6K6HAUZ9LEkLSKxPbi/rOsQkFhe/hX77mI+GDvtjW73+Mk+r3VFJq9+
YvC2DdCEAlq98R5uBvYOAI5nOvafMdQ380C45Zd2crYx5PdJJGXiSGihFmVuPuOcaLj2XfNGDiWM
QfdH0UFWG/7a/jehFROPHUE2Pn6S5z0wFvGcpWWQ9TJ+jDFEzoeHD6P3/0omdalw9A1pst/Zv3Au
uZo6HqJaJAoEidKCVHw0kENyJ5ifNxbE8kJ0M8XN3ZcJrsBIOS+91G274ZdEdpEJF40Twmwc+Q/+
1d+wSc5Lm1Oi6zfO8xvA0rErwBw4lPv81z7LZGeaOAiFR5To2u5/pmJZkLf0BA0ChRUWn8WkhGmm
tNCTIYunN/OYMZmiwrVFgZoruxfkklurTHzal/OT8ZYfzYVxMAsWZxis1Fy4iiTnJDNcNsnRgqI0
omtBpUG5bFlguJXF+eLy95AZdH66YjWzJDJOQ9VNUFGxp70UvZR1cDDTCzqlUzVWEKAajexkkEhy
zbGKTiD39QDytLikCGFfIHHgAPGKIYYWPTS4ZTJrsY4LgU8E1BTbuhr19ATNZY6wkHmdlPiAT/EC
8RTUfGfPof7Y1mcnR8NGGGrFBd/iVkrpzZ2kKoue+xdR6yNSfBHhzHNVhYP3ectquLRhdor10zbc
PpZBKLRdoMFR2nU4TgvGZEiQrhic4gZFZtn6nCiU/wxJxVGA7z4GhyonCv67uf9Gw/KjF/R8YVM3
0f+dKRXM5jieU3Ybna8OTQbynQZOo5ZFlbAY7tHNeOhIAZDW5tyeP+8SDRF34wCduMtt72s4UCQs
zf3CjB8i0A69wd+nVSnWbRJ3bYLxcnEW5IVCv3V+yjNG4WlXWHeC9w1Ui1WvP2YFlulhlXjki6vK
eE5QlB6PgSIbdsz7XFVXIuUDlqFHQ21bWrmeiDn+Ciw0bZg+zMib75xc9wsSXbgZJyPTO5WdF2zZ
Sq2yb8NqZVSf74Qv/s7N3VOt/kyJa6jZKmEmuoOfsQjsZWUbArELxG0XdO2HZO4apHC8CPBkB/k+
bKmofjA+mv5ad3svwrOwkD8tcjq0zv5gHIDIb8Sv3gHHKkDjCoRZ0pClt63Q+p2wTEsXHPMavmW7
SRrwWX97ctPlhl6REmUJxa0dHK0yLL0XwFRhJsGMpyql29xL0QT0NXEA9HcnpIIRzBm9n89ahM7l
st/m+THOgUDL1xtMuP1Ldz7qzaOi3LyIVNcUFtuzUj8MKjWg/zEy+leCzrdR/Iac1d94MZKvoX92
djUXI9z6oc4oi20r69VOBsGmZsMqqHu3appIs2oPM30YQlxJtpSUD6mhHtpAbvSR4Z5/dsHuAKZf
S8XNifHDr0tC+hnulKZ4aQLSeqlEdSnK/Vw9NwwZX9ipryjlN1sEEYjkzJ1TwjeBXoNPajTB8moG
1lP8WfOuuoZccwQ6HmSMPHZbWzQO9x+LjVXQAsnGAlC7WV86Vtv29H/twVDaJx2ucItFoTH6Sl5b
xRcXgPOzXbXItQS2E8sPr9Ljoqk+PsahAwmHXplYoO+5fZKWSX3+Bj3iLWqr//qHpzh8q/OPIAIK
1wbMtI9a7QTF6Z8Rn3Sld43UdPDg5qaa9clCFB2B7yuLuQaXw5nfuH6h0RZb+ECm1zbDJdmsqtwr
MPtAf4rOG7o2q0OwpqVvE0Qz1t5q5bAx5/STQmC4axmSngaIhdtTYIOp1GiUV0MfIR3mSvOMkUYg
WYGVmzMlSNiHWC2U5PbLlFTvOV41G9UqueCigzDR3Wv+AjVGLvP98q47p1vbauo/aqUq4RcZa13D
oLFUkFpLmjgmv2swa87toKqwO1bxNlDYvm+0DsW7CGXDIOFqi/2eoi3Zzzm5DpiF5fB0T8gdrr1t
cPZzWfidoxuIYTdncY/nG2wis61QTgxlfCg0lXWhm7/CbJ2nfJJ5p9e31Hqmr8U8E1k86FlLjpNg
6w9jEX8N0AAFeqd6RukNuY0gL5XllAsH15iy2SmjxayDJPFLPj7gNNXJkSWl9GVAbVtiRU2XPZo5
n6FMMNidmvZKP6CVwyWSPIXpgGsVDfR7vWeYUAyEd4dSJ7jSoUTxGgcDksvVdlTeMQ0Sv9ohldIf
V1Krawh3kcL32AF7yubWhLOVCW0sGs4XdlFzhjiumzFoAoiO8Dm0byDmUzM93J+ccjDxvuysa4w/
mDWeu1kI/d4gAO4pSOhZtj/sjWQyVooFq5/KrxxkAWPeMfIuuNBLEq3ZbBmoPLzfCviwWOigSkvg
PhyZLKhi5BA8WYc3Qbcq6pDRP1SwJw9TbbYcDQEzEzI4PooZ4BhgFxDBYteUXtWKGXf7Z9cKY70P
m26ty8F7wHmgDmt12hgd8O9mp6WhxO+CQNDud6tfcy9l3CgZrU+VmUSVa4N+LXAcqzNXpGL0L0lJ
myWh1yppYdFkgNw4TWP+Ee8iYviKSfInZHl+iVB9zn3hY63JDRrvnVd3EseAn2yB+NhLhnKNdEtx
FXoluOF1ZEa/y/dKifWuGsCas4Oqff8rGdGonftoLdEY98rrBz2q1jhEYk1wblh74mUP9twFKpiS
lNuDGsRy0E1IsC0sHU2kOiKz76pEOyn+Nv03gKbWpJ3pA9EHp0SVyTKsDbIs9RM6g1QmIXhi8oiP
fJBRiWBoUlKpvEGG6CmFj/X9HXH+Xvn5MAiXqpKl1SKAFroEILNIoCk9GUEa/mPukPDHccgTYmH5
FUYa2ikCQxiqVg956by3bZKnIFfqV5D674RZqDcsPEe1eisWO9YYBAUiYex9Jufxi+1/ZKtngh8g
uGVQj1U0YAjs8iOyDVRewkTaYpMCkHsk8hgfXT/w2M2bNKbMRI2QdgdrOrMzhsqdVeJVLWgxo+jh
/xcgis2qhF+dhG0Vrm5jlfHd4USAlu3+dc0hNwYyCULTDtNRLHu6IldXUv5nlYB3pB/4OXhC910W
EjctrCj+iO9mZPafQ6ixfBNuadpvuyIScQ3WjtV6yq1EAG6UfSji78+rVFfCOc0O/rY8kpnXrNNi
nfz+sIzqUhcEGb8JkWFuBBl/mCf9vk8Di/zR2zImPl3tmCB+ON7sLJaIb3cNho2q1XTHL043Zw5Y
JkSOz2lDcjzBUk7TygxQMauqxrToDCehuJ0vLpXkhZ0NDk3epl874UitzSRYDw+1tw1Ve0PXluVk
3DVNcfJ1mxM63BOmyXenA+iroRQS2RbE1E3LqUjwUXPfIpv3UijWSiZV7+EY5wrvb1ximpGCyuC9
ABQK0o7JId+mMnTEGqXW4s444ZA6TRqu+2A6ZY1OAOaDw5+gmzDMQAN/yOv5GMmqHOIYyaFLU4mc
fvDH5BtmnHGEva2jJ+wzPgTfwrWenxxnKVyJsDkU9dakTrv5wxMreDveKVZaLaVpP/Xd6J8EIlfs
D0vPmgalLarrCE5I5zEJJtPjBuZoMxhF6KgU+Lx3NoWFJbR1sb+u36BDU8ySnCrwIhGZtx4AbcPV
PX/QzRvgOkTODmySUUnWqbc1XQjlH8wiYX13/P/m8DXLLNlkHaJkBkciWt2nSdzSYQzDB6Kzb4Ra
d0SvtWgKW2/+KwoQpL4ypXMqF8f9OK377q08WJrxuqgcGYH04fB0PqAVUrJn1mZ7n4raX1eR0YJr
wfXjfsRaFJWaNXnKLDgubgt7+Pa/VOg20dxvloFcjNOaunp7J/4i8nc2xb+SdM8kZc1YESI5eEx8
cVtUf4Q5rJj0oHYKPjEHY6nW3WjvvSP5DSe4z+05LhCiUxTEn7HJT9kdZKq3CMs7NKhl28pM505V
m+A7FhVvxzY+31kv09dNmSn97LTMTbSnbcS/Ie9zLlYpgwI4PeMHexMKy1HZZBSA6vh5bijheRE5
Bpn8neQRXVri95deaOP9880Zi80Y9IiMU1CVlWLmlPIcRkcwzb+8rtgSyZqePYuS21j3h6JPum3K
F3dZRB16vKxhtX8bFa4ZmeawjSlHzU6vzPbmGgXbnE7GitdmI3+W7fj4oUXSj+c4OZUS8ZEJNE5z
k/NYUOPG8byqMoi/Z/7KeoVNpwBCeLw/0FmmLJam4GQyYFdalOfDjLfNRSaeIWDfiW7xbh59Kg6z
jx+5fNTMoK7S6AGg+ioZskL/y1q9RqJgVDscnqijJFsaUA4xylcYtXSwErBdC3bdQxCOVwkIe+p1
So8l0jgRacQJdjZNzUmm9nXoMvtxf4v4PHU8asd0r3CbsTlq/b2n30T9DvtM6V56ZamSFiKwqqRT
NpHnBwZ4uu1LqPnZn2xrULCZdW1oG+Kb+fqlxr+kVNPRc/RkTy9FE4kmpC4TnOsHYDtVv4W8E1TR
UWbGr8jyAucn/bND01Xb9UaiFqWgM3oMZbVqQUd7IuZuiNLlgIJ+hD8iSsGxdCF+STTf82AipqrD
GRpkKzX5SzLmPkryT6TnzcFpy28qSRX6tLsoBllMjXFXL8EJjOmxrauN+UG+0FZYXJ95+Cszo4We
AuLoJovVVwPssKViYOy2MYoyV4g55AC0J8Tmk/8rJI9Xa7pGeFKRhFqKS8oZrhz1WreE42ruvyCP
jHgbvYq80Sndu5wjsa19OaBlhDscgBnMLCcHrssroMBvX39LbRCAn4miUugzCWhU4VqgUK1vDMhj
WiTcnYlH+VR439Rl1RiJW0/P39XcwbEu+m0oj5WKNiiydkxCK2CUVxdvon8fzxwuTLg1V9U3nm+b
3iXeBQpZ294/r13NAL6CO3FWjqsWf2IYtdEm/aKR5QFqrZ+fVMOXNUuD3l9TvU81tP8Pyvq+MHsX
o9gE5X7I61DoWqZP2nuJjxw+aYyuOo8/lsnrCLIfVNPWvap4Tavvs8mW6NApV8fWB1akm/PM2LdG
ZngcVgxxD+LKdfULTh0fFS+5E/LTFkN3r/OtO/tMl9E+3Q0ma+ChcWfyIqh4jOmKqUdJYESvbjAb
P6qmMTkI2Kox7+brdV/KuZTn8C97jMDxrVCsQMceJgyfeTTuRFXT8EH+MYkHrJazAs3ilWQYACAw
Z94QnLgvJ1ds/c7AA8OSK6fMFzAnSlkvQR8QG5ees6acZRhfFpfudLEsttIvnj7909IEZNcrbGBx
L1dP0KeN14LuNVTYdS/WXNtKVzDfb2l3aRmrnuKQjtpeUEkOMkvriG8ToVK3bblOGxGbZG1rqc1X
5/DCJUO0HL9C5pduApZtieA5gjBOpk5nhQefj8ufyI8XEPhW7x97Bg9j9oAQ1rI+dJjBoEeJDqOx
gBG6zq03GZR/xz4wPxMgvbtvyg8ZNo4zu09yAqB/Ohl2VtUEjAabkUT+ueU7kkIYpQTCAIdaEx32
bP2wt81S6kdx/NO5pci5Lh91jPl5D+x5AIwqKyeXZtyy5YrSrBrNNpuJoIQpeS0ih30QxCLRyeWr
PNGW1ImK1tIiM858rGKjcWz3xAFLwLy47aT6vIf+TrdwpQLd+tuNvz+SdPbI4RKN1AX/b1NyNToR
Cox9avTgqvvS0hZpxVi5XjriUJ1JQHdFMPrJUNaMu+4I7p8a4JNkKdoeYTDt37baEzmUtI/xq5Kq
dfHQZZA83rOdTsuhbwAkUCsw8NiwpHK0JmMke5ET1nZ+c60Alg5unJZHG/iPkHGMF9je34Hg/KTe
TGXjZ5HZW5R8/bpYcWp+mI3SOuipPhvchrXqd1FIwY0dX2NAMKBWMldbpHGeU8ZXDDCi1tn3NEWI
tWtb3Ca08BiC4uwO7YbzfSM4lOTNSD8xBrFIoqtX5qh3moD8+31mwFPm/3PxxPv0ktybC3odZC92
4GPGR8b3y/76jzV2ggBJ0M49t8sQc++7fRxpn+JJVk0WE+MZCVBtBPfA2KCHWkMMk16HP75y6qAF
gRSefNrcipTxQaMoX0ULEFWvvyLHA04IyqLUL/iqFhW3QI/SwP2v038+05J2cR0NtEgy/8Zcu1Z/
Fs2I1iP/c+OuJFvgxBRINIn6H4GiCbZ2ljNLbr+N3Bl0B6LLhpPZ+SjRZh3jtesxBuAj/7FUWtmz
/sbhcYpew6vts0v+umtp5iwy7OEcqrIb26blNdxq0dA7vBHdsbyCSdxPzCIGggvw92965JkRVk/r
uhBWpVywUyVoSErwJlN2WnHYx+UKC/Hs3VelrxRiukUNKNP7JnpXJlenSj9QSE81QpcjhLWka+Rm
0PtSoTeESj/tj2XnnQJcwU4V+DAEn3pr8yUqDnG3ZmMTY81l7iZP3tSYH01/6bVXibWVuZFd0MlU
L2XH/zAS/xLpHnEt7UuMoF5xx9Q0qp0kLASimhnni7rOAmEU3es4fNL9P7kvK+j1AC7R19sl9U6L
E3A2WxWLBQyP6U//0gVvcjXfq9gkuefoqzTv5EpSWkpZox2R0h0qVsiUVHls84B83LMIndppbnTu
KP5gnKO+2YGgJ0HjizmjqMG1WNNEUIBavqIlPhuk+eu8o//m+hzRZaxMkB9J7zE9jxguvmpkfwIY
Xyg6nL2wgBRsQhrsGduOS2RVabXeyXXvfJDooW4R7We7WjgqhDY6ACllL8HB21BSlAIC3gvmL7w9
TEGXq1fdWRGT31w6d3lbq4l6Jsgopa0B/IQVkK0vtG/hBOestDlvv63WFjU1FksGYmMTheUpJr+P
2AY9nLy3GxSK98cFF4hr6JxaqoY13E1Ll4g6uJS5+NnN0OFa8BTAa7eZfqdVYcX7Ik4JZ5Fn8Z/c
IYFnhh5iqPKPSx8JID8oQgVI7cVxi0Vrgxdqr4X7BBBwZ/WVWfG5tJaoMoA8HQ2kAx+jM1hmv5ID
WBRI/cmjQB0mCjEhfyaH/KjNPlixDX6+gTOvIdjyw2AzIwqFRJdbHjnrhQocDaRLXMsY3aGmPjo0
zqFHEfe4S3VdKohoBuC6BgoqdllcSh/kITj2lktvANQnE9koCHM/wp//bjLWU+FnB1rZB1nQdvLR
9lcuWYIWAqm6LbyKTbxNDTXGwag1AQefzX1FehaHg2Fpe6H3751sHona0qGAjICEadSCb3szR1z7
cMbZmvUmNrG+GpdLBpCHlCRbKjG7xvoOHfj2yc3EluzCQJlAi9AsgHYbambj9RtudMXXI64ERqY6
pxpxaEjDG0bPbuFKZ78S9ipUo7SFyilp4i+EnYkclyQEVtVDDMdZtL1MEFs9P9MY8/zArfsEiayP
niHV1/mf7CgGA7q2wedFOuA0t3xHIcuthnd/2JkcqPhwtaPlxuXIBuFuW3eZHx4vgJuSa1yQLO5s
qnWFlqMOftRaK4//3ewl74n0CHzSJ6Pq6qcDveFVUQZVuVCYm3Ddcqo1IPKuAA9xihaPPZz/+7Xf
6BIsAmvT1hbJ3+Fux7QZJOiBeJ9T4mU7HGHaQvIu9NVx8lzahiKWv2BV/SGvAJxOtTfofdqxkchr
sv9rgGga5Z/d8zbFvCGieQsHWcmi55X4w++BcokjJ//ruT+o6uOYdBSPxQh/2Dzv3mxMTVvha659
hKCT3y+v9+cX8vkY9zv7rISTLXdPb3ptobWx69PRmcTqHY+Bykegi2bVVBNB4YMkDoLQzuq4ShrO
Toei0LWajyASTgZKTls+zk+PE5GaLo/tVSxF5T9Dj9aWImd/w2M9kObHkSRIP2pm0T150oqHpmLU
8CAnbOl2qxcKuQMtaUH7jQ71cPZPGKzQUITdTYTYKDVedSjp7Y/QbMIjASvdRPoBRQyG7QFUv0wi
tlRXQxUzI2DbbHWf9EtWUJFjbiIQW/CJHas1EcgNWaDsCOLwUxOL7lLMUSEPQUtdQMTPNzhJfcpS
eLtnfuHRIRJdqdkrnL/gd2S8azmbgHWO0bHYsexOsDQfGUvziRChzk4ScHg8R7YyZPNnqaLa0iwd
IDa6KVFNJ/TsmSkOlOukTwwacD3vOuSpkVDivH3TII7Gvs69UFQ1qdqjXfwlfQFSgdqp5gKu3Jb+
Dfq3makOU8eICs0lL3yTph1nVBX726GkDb8qBUFQT8TWZJxPwELp5ThM8iieBYHcxsI6D49AvmSY
T785Zskf9ToP2mVCJ+ED3wih0nl8L8udOJ6lj3JUXJloLukbSxGAGoBK4nn3IGm5OWRZ0VP88Hwc
us55dHTMlthh+d+wimvx4hQfsaW/Aq9LpjMpruyzjxkgbBN4O5UITaWA6Zn2cfL42CYfStQ/CzI1
kbWaRRXnI92+QVYBW4GaBB4A2Mse404bxmbKW2dyUmouTbTiSlb7d8QEaARLjJgBB2brrfp2lQND
S+bg3o0i65meBaWHgKE3/ASbAdbKAtidjTnpMD03VuuhBbnXq2k5u+iQCU6R4d1zho7a4iHV1UOf
PyRkUTXaBPjpm8+xedP0o7UlBOOVQMVD/j9XcFxJYoCHCan/pKZhw6YMrfCv/E2W/DGPmXG1jO4Q
zuSRGOhUqO3S+v/qDm43JV8hzo6L3eSxEts4462qrlmRnOsjE2eL8NAGIcDomPQXYTR32KWQ6IOj
WpLSzTYDm6mIxNFOIeqkyA5pXaHsjravmBE5qvSQERQR5oIFTOvaZLjMrJEIn9Ft1liX0A940o5t
Pyz1O6PIZZXy+NMb7AGl6aC5JaW0OfjbLztZFpMDUMqY3mS8BejXQnGEAqGga07cDjOpSdoGS8up
2vKlDM3SiA/OhAyOOZ77sJAvAkCezVv82v62lLJpXdkU7rODungPIx3/bl25t1/fBYMaq4kGrlXA
ojUfCAC+Asn0ihpadgXr/Qut4JAUdovr4zJQEeIeyU3LYQ/7Nwi/2JV/7xXCaJCn6dp+QvDcZkZ7
W1NmnzJMdr2GfP03d7WWNvajZ3SUDGEQ/v11IdYePbxwO6feIDNLpqskEGvfSsRsFVfMv5Q01NoX
55ERzImFEQAv2AfziNrRJO7tnqKnkS9M4b+fILnNCaiMiJ+I/XZ4ButqeUabYWHEzXIBNDzf1flX
gYUn+BHS1rNCCTuM0UO9MX89GYMdVkFrZGrdTpnHOOnL/pbQKZxTU7twn2rqez2wUXgjkMW76Fd7
HbWvEtrAuc/luzluQgm65bZSNXp8VGmhxiNebLpHzOmLSnfF67ubJhJWXBHxSpW8BWsYptVRfX/V
FWbKux6S5hJWJA03wfE/j5AuaitO/62j4UnUNHgfe1Yh8enNC6SjFbpfbfLcdNE5wOdWw2cIoHz/
pbqo4lVq6EpgcbsVaD9yzPss0HwR52rANbCfidaJCC1pwUSp0aQvMSwIV/s/acUk+EzOniC1PrSv
FQiaoLEt3Dz+epFidmCaMozPYk1KHAES4ZCJWqQ/r9O1fBoh131M8CjdLNtyf2ZZjaxu3ojkdiF9
qn9gm8cF4f4Hl6ECOMvuWvkkVbhHb0hNY02U/Iw1OzbTZEKiWPuTz9V2GAu5e5UZij+syCOR8AN9
GRv4EYNxrLN+Wz5P2uJmf+ZtTjuaM6laH6c06RoxZLZk1LSeziekbDTAHBaVZSpngGGrjNllEr+x
DiSNjzP9hdBqmxN1zCwj25W1WRlFlOHYvW+2qaq+AJyUud0D5hi0eNCICCdd9vpcLj06FnHnxuZ6
7xlMo/3ZrAG83aoglG/prM+GQ6Zh82exsUYE+I8xF90uyiazZcEm57VLstYVdP82lFCa+HdOz7pl
H2A+J/QgDQS9UpHWU0RbmEpvBniuNgHwG9N/PwiBmt0Jdvo9n55X1KMAO+XXnfvr3b6NX8GZITce
hsy7KoVos1ZjxzaDsc7Lzp+9x82kZSqJTmUhgH2gLg2DMZEKmuWdm4/u6MV4LG3SfbnIMDhtj8yo
d7jzHbmhWIiwpJHgXgODbHVtkFZPZ+y3X7CYBdfnXA1YZLhGbauFFQqTSKj9tK063lSav86HRt7S
uuP5VqYLUwzPkEgarc5+VNNQuaYtdoBUPHYTnCSBa2Dnz5RvgA+5TxHOQod9kfb0xdMa5HfpUu6L
eqUsl4XeMyFgeSn0JCdIvEA9NlgW0pI6GYXRCwHzKlzbcSwyOukZku3l45pxeW3tc/49MISG80K8
G8pDgI3cpu73ESyB9doW5PU3wxy/S5jG5vkJ4Q317Zt2WZxjz08zSEYIbOPfG5LLMFzpDLz89uwV
WcQ9ccyG3fdWZqczp9h6vOemY79dPWFgHSEr05N4kenq1fZo/jdi6yoHyT/cgVLYacCRXVy7aKGR
FOuOLnN2lrglPqzdeMxmA7XhUBlwha34HQO/KUg26RAMnWu1Jj30KwPp/tU+6HxAEpy7zcqt6EHW
kinhVFBKu1Gi8p63+riy0SpH8XFhHGVlsNOU1rK55U70fhVDStITtlMRn8w/ayi1l0+hPGSRBSfV
0rgV/HYKci786WW3b3LU9sxHqaK96dqMBPwpDO92iIeBU4Ihl+e+XQu9MMAiqq+596RmiWGCK6tV
tqFs8SoDJycZ0gdinEfHWSuSb2CWi+WSoPWWYKzZVcARv9xva33qgUKQ3CvGjMJGb13B+Nyr3pEC
83LPzBVdY+3zwx/eqWjdSUygre4yqbDT056nHbjsoIp/3yj856aCkuUkze47geZHaMQxJqB00z91
X+8ris/XHR7jPehf+M/BPZyeaKtSXPRUj738r7t4OJUbhc+c0yiSUrOrNeXTp6OpHEL/cI/d5MlV
Mobaoh8rYOztyJwjWozgyZXMzdD/SBEsSC3pVAm2do4/LpbouDRTJkI3OAIytbeUj+Zy9m7F8UKD
EX+p5UOqXnwqcVqR5cBN6iQ2AIj51ex5+W6VD7i3aQHDJyGFonVFUt7oN0pYChEO5ogm25Bth7vu
OV5GxPXk3X4UocpiqneHv2r/9tPXwm0BVfujtp8qbhl8EbCB0n7P0T/F6OGZu1N3CcOXhAmeb45a
qrHuNlc3fz5i4HlvzWUYljLxa2hsjB2lNR/KJA0lybIzOi5eX1eVprmo6+W3KC+zeotP15EihpDo
VcAKqQNJi6pui3AUe/S9GNS4pVGyAreUM2sHOKUugozVGjo9Nu7to5EqnVjqSzqmfHux4y5xz7IK
PrKh8qkW7YV5/Gj02mWRpmz2W9Jp8I5r0ajcantafYsT2XIwcFWRJmK0VfZhHXcnCwZbaPf62RpP
F38LxHWfockugqipnXQHWrt/zsXEhIcNxYqyYw2r3DVI4d9xcNBJj/9KIBKxOyc6R/Inii7E+DXk
LWlD59+rtxd+kU+7G9pnRZoTp9QJH0cONsYIGQAw53Ve36d61ZdvGcGtR7DPtOnnELxe9/7/be2a
MEL9dosp0wCeKlHSOlcuZs+FIPvAchafwNtjNf87JkGzg9xnCtqE6SA1CyCIN+WOGfrQhsdIzNmh
O3vHVv9dZdcRxHrHgAO0OYhvA7qZO1Bjvdbc8StfD9kTx/9qGIy5DSs59eB+rRwpUZ//u+nopePc
47c5dEjl4TYuk2iXsGEmkQBBE6oXLX4BlZZ6i7bAi2Vo9l78NHiLCdgCy1mIF/p0dOH3L4VZus4E
TRHj3rJKUf0VkKVK2Ivx3mWcsHgpthIm3vSKf4XKSbHOSW9wEcqlxROmkJPYHuq1a7BamqWVcIpR
5zyCQHJbGpMy8wD848aXqLUVRN3JLYXhIRzMjVIgqkodY6moFbXnQwY+vxIM7qS5zKqVscS48BbT
llK9cB8Db8CfFdP5CVgu+Z3j5yJqOplfbvobDokkSPupeh4BGLH/pZDNnECOLeU+nP/5JQV2aiTy
1zkD81CR33Pb1Pnbi5AJGyCFnGOeel4+MmJNzlHzIcQk8ikr79zI74PUoO8wKJJLnbfY/Q/NBYS3
XY4lWIM0mucFNN06+1nztjJwrabATkNO032r9q4ocUCQnk6o5fPAo/1ue+pBu/XE7QC6kpL8FSqI
CLXhlhaDx3Qcpyy3p11tHrndXG49SdeFpEQbP/ErczbOZ2wjUQnLYypO0xZJnkZURCbABOm6OU1t
Q4p2/EauTe06wN4+rDsE2/1f2peOCCgLoappQKUo+GCMkELAAu5Wj3rARvK1EovPMPYGdHt+9gya
qLy/v1ImcyrqFupFw+/qJ9d7koWqlsQ2dvDsIJ9wi+hseCa9GN8h3Iz13sCZyM7qbKlqsOg1yBqN
fs00E34dti0sXSr+9/1xBJtI/o0XwQtiTdIXWgQlrwUtw8Aj6wTG72vF+An1Ucw/ax+1k+v9S7Qc
4DwvBnZZzPbm4SAru1BTVBrx6fq2hfwUE4Bi4cARgUb3Jtmh9ennf2Vje/u9C+xMBKLe2xuuq9dc
W9xVdENk26kYHJlH6m3tVswUI8FWmzlU6QNYWRfhzT9+LPTVu0FJgXhJPBEwB3K68JwnBH2YtPZS
1xHp6JPUo9EA1GxFXa4jDCnvrig95Yq7z9uPOMzEVBnEaEo5yH9eJJXt38YGcWprzmeVXUw1XtSM
lCGzmog1M7JKWNbJ/LPtsa2vbYYc1MrWzegm0NwVcMI7TBngXtHt1B1/h0cVokm85DTKh9Xp6bfB
AuTebZWKeTPgBrz/qb6Fch59oh2fZAWIV4A+NqzXCkpBCquDOKCOfDVoWh1+ltJmXP6e2WRRreDT
ToM5erLpQcpAP2g7Sc0bJIC9w+IgiiP/3gvaCTQhrtEK8hBRy8LyvYTHCOlHMeHY53VMIa6DFg1a
leSuDnBNLWdv5tDI4Cp0wNf5aEYr3IKKa4PFiZKAfCE6hnQm93mIN1e7rUnMVVLTdM7H+JqMWWVF
W5u/0zNeQz8skbi+RN3vY3acRNrnS3CemAultpU4qc2KfzamUtk7JLgyZF0KjHU0MBtJ1JGZpBfb
i5e/juN6scr5ppzjOQqeCKqW7CyZt5S8oGbeDTHnY7jtiDcCgDW4SJbqSTomywT3sIgrAh7oWBxc
cVOPeQP9ozAESMgCfE9uexNNOkZwl1fcBqrkAGWB+P3FRAHsFLBdoddFXSoc8Hqin5cYUrk1siDC
X47PBrPXEHBAQ2jMu8/flP4AOvTa7TWP94dxDQhqHaY+PVqL6KEzpPlZEdPyZLrd+vb7AzaSnehx
8vhVAwbeDAFsXnZkaR4zEI0My7Tnxpo4yGGIjhoW3MVULya6XTVwbEIJO8KK6kawUV5UNhNkqpAG
oXTSJLBohH+r7UAWVCtGgGAOlC3vwPmCIv/K6lL8f1ug1gOYv7xEQ4wp+Y8KbkqrUqGRlTYZ+ZiT
E9tsFHnc1S7SozikXMcHto49puWde3NooN1Q3TmQdG4ClsctyeB9Ak0GS1beLnv9dzeqqE4HS0k2
dY85c3U9oLZNthgEPExAJD9+X79BNg0Zw5Az5BQ7q8jB7FrF100zzv1rKi02PQUBP4cj5r815xWh
NKGmNs1RP9Is3WE6vy5qA6tiNVJmrPJo7ja0+AqLWVHwFKIeFmovR2htZP50jPuaEe7ghmti8Dbf
RHHkyz0tNS32g72rOQqdZ4rfm9RraBuBeU9yNapSIr/YQvg2YEugQRqp7LIaCF8UCucLuoybyKVE
yPCc8kZ7DXPlUJXc+WRqDbJVtfuf+HdoZBlPq5IIkmvpPfxTePJk7Sj+u2L3SdmAGMuaha3JMx57
HIAwEUPzISLafMErXpZWcacQXBRIAqHC5bIfzru8HHglftkAksr6/mB/obo1KQeW7iJR23zxkyq+
Yu+kvIPew4xKoEnm+qpmMGnQ45woimuKloxXi7k82XoDNLY65oUQ85BIYeeASt5hTdchTSZ1X38p
3RrH81mUTbqluuQGVXQXYGxkyQO+eWopPXkPUCZoopKe6ZySIzZgT4uQctbvhe9UkEHRX8TrEzeh
Ns1ghYhNSFKH+RE+fVuF6JSk4UqHTrDyM0fkTMn759felBCNVelQGQbswyNkLIY4RGQAtT3hE6OI
TB0JIWX7iZt3DyrIjknEXZ49epSBnEjGkhekvjij7tLdM0/HynaLM/vdKEofQS4qinjf3QVpN26y
FgUiPqLQs+lAQ+FKZdqqnFsqTuLZAe0eg6CHq51PqmxuouLJaBTB7IjhPPlcMOUnjVwYxKS2yMkn
G1AVP537Vlv5cLsuAJT+dZJ+Kds//s27BB9do/tKjvDkry2IJFN3Ku7XIUbhkhIdCyu2rY3PrQRF
EcbD54ZrOkiK4YlX2f1O1iDIIXhgM8kwctzW92RAQ0q0D3zPhXtg9Vou5vlRBe80Tm2cv7rIxiu3
e9X5HminEW9IGZUM8cPIvNHUubaEsowNJU0Y7csqOef17NraH5tRUBl7wEGnHroAobOhX2R6lyf2
/DuikG6APOI0Y6wzeHnG6+oD6Wc3ciOOuG0d+E1Gka+4z+PuEIln3JRVHDqXUymiVS7M2h+kYPt3
sZmsYY8Vyu+d/JN0YUKLqy6iiVdxQvxMmrs+gbLtGFSY9yiO43AwW11IL6Q153lZbSyXjk0ZQuY6
xCamLNnpsxJM1eqA7Qx6IQtqTF050jmRb/dqywP9QKLto679zQglIa23UvxmuP9ZpQmGfTeK16mo
3fMvqF/S63eygFgtFTCi1kkWC8fZz0J3QxXbZTwR8Qi5rSwyfRJUK4QTv0zIV8K7Sdr5NPPUDAiN
oit32qmIVk1zE1sgK3Sf39i3XfT1hlggLtmbXxXPBauy987H7PIWTdAeFlVyZkHla3ke5YSBMbi+
O53bByLkl5WOTJQL7T0B2CvCwhm835K2sZEasD1spU0mSgzGOc+2paBwgPPv4Lftrhf+qda17TJf
yC4uZ18KDlt9wtPyZW0rd2mhq58/n5AxiURxTtNlFyoHA7uuz45YV1aNf2PdyRvLV6nwN4AHd8Pv
fxonbGz3Uh2dYVsN5rw0U+2UJOK+h9nVykcsU2H2u1ep3OjILUXgdCRfL/mraDeRZ53uIZWzwo2E
qt8IuYDlDqETJ/GRYfv8LWqVbNz/ydZM9YRKos8DctfVhSYI5yByzzXAi1uRrc/EmnCjPqHGgujZ
58qR8ginwJYgPIM31YB43koJmh+k9oJ4GEBYMGVjg6VpZkFGOz+3LbvIaOfV5LJnlduEnyRy/LO7
ldJyT6ute7g+P+WVP3IcNmPqlxOR2YjZOBt/eil83oFX3FTdozSGUnNbFTlp2immWam5EZjrIzoK
MLlpPdFNUKWfb6RNaiBy/t2uuo7rHh7R9rlId7YlbrwBgByDBGRWCaIZ5boeqHyXaZcH7lA43/bE
TfGvvqgFjhgPrmDOldjzLTJp6MGtvVL9R45mqyH7PYnkFGlgzMVsgEVACWFp9aLkT9V4W1u9mM9p
nAYHMdNelLS8uW1FKVHxgzyPP0dWojxQ5fmIQFgd9EhrZFiPxtlTbQiVZwvjaJiXpFA+1LfcCycS
i0XBiJtrc8p4YBGIPijuR9n+CjyIyhtGyA/kw8Vzni/dKokkc2J9qHHk5k/2UKp6Y9kRkKGXpLa1
Ub+ydL4ogPbjKMjZUtMcGv7Sj4a678ej9zzDxwnS44sJjsPV9wDB7w7RTK54bg+fEhQnLPU0nF/o
f9FriDWPIPFTnRjG+YD3rmtrHv0S6XkbPccjV6J6Co+JS/+I6/R64cxzzfEFNlCKizuUSAHnZqVX
2IKGbCgxakBPhgFpi9+Qlw9RgPb6sUbHoDIA3m5egcZAiuYYbwNwS9vkoKwTVBpiscGagJ2mm5jT
5sX6+Zw1hdfAR6N/PTyTUyUM8e2art0HqxhGSIxqGexXuXkrJVkc8rGoMS2MOgJdMujcmByC17yf
W0qgWNBGLXNSsLp96SLVV3hO8Sfwb+yv/5nD4yiN6qfjANKq+YdsGrXWSp3N/nmpZmpn8IwqoMYQ
Vcj+hIX3CJ1/pcs7RMxhPMJpHXC5a0mkq8J/IICB6zaxf16ZwI9V082JHxq3QfRqLvQgGMkrJkyQ
LyDFoL6xH+JsrRMxGBMLm6Sd0312+QpjWsCwdNi7kqMT983W3mdf7d8lzEfVBMsGy3fO6QkSvr9o
5LgqgvDei3wnRepUhYQaOxMA1xzJefDuB9jlfy+8XiMfir9r9y8EpdpF3j36Vnv8O353pcG54n47
3QYm9Yfgwp5wBrr/hCC8QeVVz4MJIkJk83q1gUCx30k6ASI6Rj2Xn5L3gQhcj636xxwSsbITe0C/
9b7mOIc1p08yTkHp04jmSCkjzvIu7K4XCh2UXgn5graYQItQ2xD9QOQFhPhqC7UqtzHgpY2W5/9P
+T5Fy9OK38s/U44fV2pwu7MYroaXVwoNh9yf7DDNJgka6KpbsvpqYyOOBDAAJjT8NlmADFp5GFci
RkQrdwHe1KA0/+zC4v/aSKf5QwsPUAjgwOlELri62QwiEIIT/+4UKjISpU5xZHklRIhaQLkbqh7y
o5GktyXRbmLKhZ51UG+Yj73Ip1HR2lGomVsRPcZeB32vEp/PYlyTw17TVsSHbUpdIH2X3p8nyc6A
dj60sLdVze5T79KPKPSz9m9FqdnIjOpDTqcSRvJ7oHct00c8o6Q9gmJqu4A7qWHDCfK5WWa1aEg4
9kB9GwWC6clC7kxFUc2I7AK583mV1MQ8Pd6R2euq5PEWUvtjy4V6YEXuYBle10nc7KhVW867DSfL
GN06FPodFKtfwUb/Jy8rnw48TVOlfJkccKsPixWNooV8vkl3zP24fCfynOUMKjgHK2fKVtWmR51m
5rstklbcwz1r+vRnm1eA8TeYZ/S/gE6329ZN/fpErw30T/NkCgZ5PieUnG44dSvPhjN++t/CnCwB
RoQIHE8imwnC9qENHn9/drM4m91Si5WXrD6O9bqBJh3utA4rIOem2IYTcKWumcvNUEvoS5Ev2Xoc
So1Qj10HMwm46B3uuxD39fO2Z0RojJEg6XxaftBaSuMmCblS71EuDZx8XZxvOpDhISkQNXd5Q+g6
+jOjQ778vKll1ZGvxT+pLmPo/jihfB1HKgdcGRtv8BDDPEuiGB05wjp7CsJudvvEtHALypnsR2hj
/hPOm+jXRPVWxf/tYwME6u9ijnGV9Gn9VzOpYkvZgaZVyCHuQUWTmEEbQ8H+TdUnqzJasXUtRwkk
3QhQ/Om6QuLHoYWwvf/G2SWXcgCxh0dzsO/2ikt6BXJs5r5upcGOb2KaGDQ3LqoRBVWQamvOMsuK
DnkL1Wod1grVd0SnNjc8Z9fn83ZmPVKh1+czjm+ynkM57bKXfzoCD1TYd0oc5+VCHHrZVJc4Ptcq
WEUNTEM14AHINTdzeC6LQdqo8IfHHLPYwiQIeMK/vnX6gZAWsy+gbkhtf3V1JM5fn68IJI7GXOFJ
6jBSsIt+cBeuuK5P7Pd7co3GrJXsrjUVDBIzgTeDEA74EHi3pNQoymYShU/IorkOBk+dO+dIC84K
SFkxcZfj+lyzjDKBZKLLBJtjtBEqf+0AbXJupQ0oIHSrZQSGZPtvJaEJLxzqjLa9QHmXJFOXEeA0
5/GZU+Jq5E2xrVZHi346rzrbzY+FNpzVCUFzysuWzXo0v5tbWsgTFMbRMfSSNyCskfD6rmSqmvks
e/41yLns6dfned8GoQjPxoq3EvPJISDwSV1uplIJFHoRNFRCuQlCRfzTUU7HUJ0QakMOUXO/ubht
Jo28Rl2xtWxp6UVhfTK2wIIPAFY62f/gwNdjHOMENmZ+MRYCgksGy2KWlufY0OLGjkUfS6wEBhZn
mR8trQgMsHci1fi5A9tZYyBfjesi4TAQ519tcuj56oy7NLnAkT9Y9bK1nQBr61EKM2n5fyVcZvQZ
JJqGGCQ5jy6KzMxmCEymHg1OdZU1gBizVQoroW5jiGBDBJiEAAZ7lsr2fOcW+EmvHScvafrt3Blp
WL2RZVCVRYLbSAAE6Hj91mHXgMNSR+t7wtRvO94RwiDWh/EK3f9YJUrrkot0w+f/QAe84uVxeyat
Y/gaMYqn8/blNmZY10fDLO+YIWY31mwCwbzlWD8wVLE9H/khid8ryf7D5vt2sp+J6o7D86W0k21d
i8Q5i9qRw+4wzVGVulFboliA9rCKhsWh4sv4gcYKWDGzFiI91vY2hL4wfmL5ryDZW/X2suH3xFWG
2fihRqaq42H5f/Bxn79juloATTOeq4J5csMiMXthUnZw0O/N9S3RDZS4scOxG1vpqY+INQKvHnZ2
YLJjFKtB3jPlgjAknit4dRbFB/Ij5uSDDVjQuS2g2MeUPPpckHeiZcSt7XvbUMyea1frXqA7AkA+
QWXW+1+lSW78UawWnlK+4J0NG+3i8YL/dTsFnhEWvhWkXdVS5pRPddFbC0TdCToHwNfni1TvuCbz
8BliT6MH5L28KHoteB5JjVwKmKLkiIEHgzcCbEty8fuWcf5VOdU/xMh5dsrJKFHzoXxX4cFuEtjy
gBTiRR1rLVtWwZTWqtlF+Q87vhTfOp/zEyLXYfLR9XQ2OTkglscrBlZCEaPWiUWdBQb2lwiROPUf
04Vi3ubokv9YpKGlkzebJWQ/cPwB63tmRdhuwrt35jrBNibm5eGvY/46pP/fOwL2Zt2t3mWx2pO4
DZrRzrfAbYW6nRtpyTKgZlgeanLZqOcIGRldLqyxCPC/opMoY8CFg3T75zO5e23N+nHkEMfRxqnp
ipBBtcfNaT1FjicfP2nFkhoRnVO3CAM7nB3IQok8Rawtgtktqnqv2NdZcua83LgA/vFucYplJtub
GAFM8kalJTCzlcS+h3g9AFCZNeCoCXhx+QlyE43tbG4rcjqZJNUAPAkT1QPjPQmlET8goqi1Kg/c
VktkKlGCysw9dmUMHDAwWe1r/Shskk0v99TUbY8V6rhA89ZI3a/IQ4MACN+mnXov9K5AWUKZeEmg
OGnkBlws2kcV4u2l7aB0Y+qLTGkvTGpbrG/OfakVkI6FCaKBmCUbFkNRHDr8o4PNaIgIE2ugPL3w
Phwo029+PWOMIEA1cK9hRl/Vw26Sg8PxOos4anLdqfmtrvXEzsfd1LhQxH4DcknvpLkYnUGnB0Ob
JVLbp895O6EgZ7jBnDYRVg30Ud5YZEbCuAl2gxr4FEdxKVjZ/QA54bvEpeqGuiTXepPR9QrDYPY4
gteDoenIOjuGW968wBkbnxCpheCViu2irKb6V6q1jXnzIvn046TIz0s3ipGSLAWLMA21R3XRG259
iQb3bxuDiwobgF99AnYd7ctiH3+onhBZRvv2oNoB0ImJD7Qq1ynZaLsork9VVOlo7tEGRnlDkEVI
BnQLt5x33U3G/t2MqhsE5vH6OH2JmEqpqByLXQTsiJm5GMJgS4VjtQRC1HmDM6fi01kcVP5yg6Sm
d9xkSmrLft44/gBKm8ijaXgyGd1jisNbjMV6AGad2zQBwt/HtTYol6w96DCIlwJDIqjRG7G6lyf1
3zIzn80ihsCNxbkxjuFEJkbEef2mzr3f5BYiVAMBy1grhqZxeBcAOu0yaB+OdtE9VXB55UhAXLfu
ME+Ixf2PRiv2Nj9rzPCHBsGDhQtPHxzNBUecqVvaXyivzgx73a9XVdLVIQ5Pf4VPPsY62qdZh0L4
1IFYot/Pc50GGMkqPep/JqBJi+Ir9BzM8LF0JPrwH3YVAOGbaPD7GeaqPwe7xQZFU0MufmkX8laY
5gljFWKxmRG/UTKqErI+k+Lqz0tDtKypl5knSHqwUEBFR4xr5s48x+MuxyDtCMqHnsDDqVjmwqjC
s+iVzdxc/gIexAr+aedhUrlbzpVGye2eHXssEF1HldRLLJucva7Az1ZvjMgers1/ZSrt5lU2q0mz
q0MasKYRzos5/P8Sprl4k/rCd04Paxr7h2m11BSx7iW1Wof3DXwmprwLyjxD/bvY6Kl+rCv1rDdF
hsGTtoYXKjwDaiAXun5Ji2yHtlI80wF87WPBuUPz3PoyfBaW8Gnt9+2UHD3BFGYeWZFKO786osgc
wU7oEklxVteoWgFB3vTHUv5ioRF3i/Mx6TBhB3ZSh1YBpTVumk3tI1gvnZsGMfxgC0rR6IfA4VrM
s2LIKL6Jd9RkDKRXI0rARNA8r61QymnGVfvknOhvO/gyMTZcirDJvoy33mr7oMoQTE+ZlpJcCJ8P
QVe557seg4kDA7oUtBkXXlbzMHvE79oRdLckae4ebRqPW2lqeVCFgBMEdSABAb3glgU8przikaT1
tUO444PkV561B5eAPVlwSgyonf8gcSGnUUHHkGC0SiyJwTwiQMJYg4AvDZXpLESbB2MgST1ZZ9OQ
8gSiCUcsNMcYpdZsW+SsxIYwolWxyWe1Y+8W+EukIWQN06bnOCUOUHl6qZsRsb5WwLk5+npBJiV9
Cz2wfBYCRKROqjsbpu5WMX4NX/ujlhWkp0XowpXvfSmhRu58thkU2EDA4RAid5viN+w3Ctao1V9K
UEHTyOkwgTHadC8nED2c0UYB5Oqmj8ZdAYXLR2Vj42bXshLhly/ZgixtEJs4NYHXKndVndeF7CjD
QyYs8u2EP0GlLUbPoMOnPmVg4dgOhtlRFB1gQjfwh5fO0DXK26t0158Wc+DVq2CHXaVMc/1n/xSf
6dNHmNgrViHVS+qHdbn+acxFO8+umlbY56/PdonycNZepCl2j4ehLplo9yV+mZb7Xd9q0BVfhI8k
YINwEY16RXA+60+E4zy5PP1QxXb11J2enlf85jEJs/NqUAMkVIRIHra3TsA23xIo9qS9Egp2Z9cs
P1rjETlivodgTSw2eVVxx1DiGlNfvibuwRRN2nmkqX3/CCbav7WWxryzoEQ3GOh/HdUx0sbsPe5X
/iCyrQa17K3IYM1ZR32DejvacvymoqLSpedi9r9wcS8XaJeNz1zY84jq0fMJ1N/9Ip0rZNoREmYE
gIqsD63VTjuHwvLHjdlWBFOJrOWldrn0lbW0H+R+nR9grdoGhTNJ8b4jh9HBZXtxoWa59S8KQTU+
K0J4AN33d50viMhkAf9RpkoqKKHa8XXFXacROu0uOWDDx9SjhSYMMgB9xKAr/a9BseR2BvgCD8uG
x1DAk29Uer3fZA+R7lL1++DaVgRqfxeey1g0g6CH4nr3wHulfm1qeewdTJTCzLVZFKTQPPYAVr+I
dfdTIpLp6LFrrXMnK6ZhO0LnlsyDdwIveL7FocwKfELVLflSi3j2QbkvNSjaGCzF+Q4NUYzAS4RE
M6NDJSW2IFxSHP7auJ1QKFOHhDu6shRNIXSB9DXVwxb4fRaV6vwGqHr7xKahQyC5cCZTj4fMSS/g
kDRl8/+zarXRX5VRHHymrz53RLqrzYWPoiY5hRyDxBiaj2EDD5giQ6EMGJumCxjxCBdysRMh/OX1
13B33xWBKw8l2Y68L3W9Ecut0ACjEmPeW7FolbfU8kfe+iCfK4RA8W0eweBueucPAhZ/9CepFelS
vYi2MLHNyzgLExHTSO8xHHriRsVn3njCtiT1FiRRGI7jKDImy1dDfpTYeyVa6+rG8HFSTQF6nnpj
fnVB+mKRL8uvSoWnzm7b84WB+rb3LzBZh7hwnrsmeBDBgweX38smftjTegE4zIBoj0KKjRfHBBUB
t01EhnWYQXYP9eZP+03732bo+xKgFodLBooP6BSvXy+3UbRltZtdC4i+l97fgVgBq8w4nFID5HFe
/LEle9rVgEgudxs5h8Zmb6PDS16u+NPC+9xqYDF1aUu3nT+ZC2b526aOG0ZGOUFJqLLIAmciwjvb
R1PrxifSN6giAyyjnGDEeWZqMIqy61MCHFIKzRPfoR08tUmY706ynv/DiJvMOPQxjxbI43Tws4VB
LbWjC61exbd/lziQJ+BzecePslv+AukrUpt+SR5Ge5cZxIk7OFX/QhKQVjAyfwG8jkNvmLWs2j3b
P7ieOu5nSP9zDty5Zicg7zj2Sh41fFQ69tgKbYH7YvbBLXeU4XpMHKrsVFn1+XMA4PF2lIChmc2t
FAXKOOE4OXS7TviAyad9A4kj64k/S31zIqYrW7jD32JqdeQrqr5QqY1B1rUBIaRD+HAHfdakYMKR
gWv4ZfqoJ3gQ7FyA+KvJy/EtXmcwR6mEwN2JsdY5O813+wHvIRHr9mAoyELVpUk+JCppj5QEAo8g
VNoCNrjJ+fdW8C14IRsUp6YVttouDTPSxNZu/ytkJJCRlRdeWJFL9ztlRPPc1rv0XF9SHWxMZtol
FIPFTrVE5HUlbyu0wh06zn7ldRp/yHZX6zjFpag88iriljxEG9G5KW5wa47s6iCq+CndY1qxG53s
icjUM7z0kLp0I6x0KZ1VWejShGDwDQO6bWxQ5loZfljmcg69ejKB3oyJBP+5RC5S4UqPAJOMJE5O
R20mN267XKOBV1gtGeXZwxnogVbfliQxhWqcOfi5RBZIYSkockiN4IiHxR1jvyug9i9reQC6JgDi
3zv6+GQX5xOUn80/1SA2YjOijjIKOFymEotqL5XeahDe902c1ostojYUt7JGEtBkC+ATWqJmrKM8
RpmM2pyr+cGETj7E4Strf641tYtLUqiMx0VUzBaTVID6noPNCuQjUsVbYPTSRb45RinKXEvPMB1w
nSSHfeTNDAQD05cAaWmvb83uLCTWe24sdhT0VM0GZOXgJ4ZWWkmJulOIYwdgXUSV0BwARBaTDEtD
VrdE2Sm3HUhIV0EhZVlv/KqcFaehaJ7I/iHlTEtI+v9zNsOLsuKYpCpYzliW3Pl7ay/4uyRZPMCD
pDT/VUoFj9kYFw4Es0YRgBOoMUh8rrtaLYkCNWaEXOTIYTOto8kqoJ94Wo2NPvkv/g2ExY8ZCJ8c
lk1veBQjp/SxtWD3e1v4adzCaSuT/Ra2UTPRyV4LM5IKSqxo5PvPwICuunV7jT7Ys8PyHzEZW0m2
vbd+saSv+3mKZEGaIdZcrroS5+qYY+TtIP3MkPr2XmUrCTsWAwrlpZI6sDB8JcCsJZmCt2on1jfb
liFj7Z3ASx7FD6nnEFoQ5ha61EHgYfmF9jUMtaCX0tclkRkB7jTAa0w84xnYyZRDTVhLkr1buCP7
EwBO/1YOb0L1X/HcV6C4yZxzA78DHDlEITbjmhVbmS3K/F5MeFt9GBGztn4MOA0ote67mqeSecZh
houZITGrIh9RALswlVsIZUgW1ZrJTw01lKo86Qy718sZnCaHAkqWAYb+YudC4DZVMXZRuZwTqwUO
AY0lD7Qqnpe9Tcr8MpJcUo5dY/cINshYugYphYJSlb5uNuibKmzmtlCUA9+2QysRioP2wQJlfSBA
RWIuKCnTystTFGELzTEPrRn9R1C+xivp/F/qse4XEkH+dzqKm2qfIH4SZ+CK68Hwzx7LrPmm2jx0
yyOqEoROsuD7y7f+v+X29Dbll73cIcI1tV57WDwpDbFZyKUR0/VFw12JQsCZiNj0FpagmGOYnhSA
ZY5koBDUR3Vm9OLmOMof3xxlEavmqtSQGKt6KnyPAyqEXJNybBE2WFJHtxsa020GI/nooXAD2Vl6
iJHPKUmkfwPSw4GwwJOYxUKfxcKsPKcvIHZ0VuYwelpiZiWJ3yqej/m9LM1xrDh2Phq8JFbGTOrq
JHe22mBjmlUO65N4tQ4UF4pVSshNE4mE5eg2V7BsDEfOuIGwjNAaD3VjKYlCQbkIy5Wq3N9WUZwY
HFBhYoMAXncjYuGh9j2gS2BGGhak9VSUKogDnjzUXdm7awQjOzdYNerEA93GxNbigW5m+UAaJS8O
IIdqgVuxvIVoiKJ32rChxqZTq+SzP4Cvk8eruq1y0J3fAdZDTKTVvSqd7VhtA19RJqJk1poQVT62
6MsCaSuta8+9N2wZaHdLo2vdMytlNjEwVkFGbY9jayA+rG348tLL5xhYZ5osJkLRr/iKhZ9f96FL
aH2sFAkU6UTop4eYL1FpqlFGQ4+6VJkYw40g963pX6aXio8YUkXC/WklpAME9eYI30v9hmDjyCZj
OMhbmlIPIN0tpE5C4IysaWdgV2FOSCitsXeuPoWmnynhtIVP0jpgZhruEcZJFyf1BRTuZrYZUSi4
SPAIiYsu4tfhy4HbDRtHcIKU5f9I5AFSKOD4NDKXdSptMcmixWcxbFl4DSWP4sJA/XBSmUF5s0yY
CGpL6j5bTc5ms6m94bezpaKuCPIU3Q5NVNR/aIkrZU+vZCnhKk3dW5x2jjzNhIQ9PUUGhJvjUW3K
5brJtSlnCRaaBZphjLDEFuJGIRwUH4sphwA5uXdf2eeU4sk6wAXmz1NgnWAle/5//x1++qj58lLk
alvtuIqpuMZgVwVzm1jrkb6M3cL9753doWMCuQ6DhtKWnCW7ePS6oUcHq8cmENrV27zK2c+A/ijp
R60mRbuvEtkYNJZBrbw5yTox8HrCt1YXGRltjRWb/7dmxpJAbzCqrX2WuM1eOEYMNeuloXHiQvzc
x4T3A4RGdDxtAv549Qf6ln08czeukIXPPG5zolcWY36mFdAWtVVWvUesP5l2fKFFi3bGdst3mLi6
yG2B80aJAclNR5KOcjFjzUmpU3/LOtvAbG4MglnRzno7B75JqYpO3KF+31qRshQix6lb/l/WMmEn
Qx0Gzj6eVwEvr096bTAlymAhya63QcHq6Vq/AR43met8D+9tIJFKZW1iBaUZfdcP0SCCfwDYT05m
sCHmnvNxPicpO8wbZ8edABxkSqzsVklkv9Xko330UCUcnef90Fx+hGlDj+GkXI78zx4fUGIQxYsP
XcGrUv7NmssqP7kNePg4CkPQwfmrnivxaH9AbwXQ68w2pQtlIYDYif8dK80/tM5iY+zSHipl/m5h
KeWzQEefq219B3oyO2Pf4mUSQzZpBCGX/Ha15qBV121gZzMt86xF3aLlBBR4IjGtPaZUk8+eDtwq
EVnVrY3GBbm0dZX7Ak82d9F52BANckEWxdI6mtvIieJ4HURwAu0pDJdc3/DmjfFD45xtc2xBbIlb
H5iFmKEuK/+yORO20R3OPRqNiNZxmogwmlDw8Ughfi1VnnQBtg/mJWSBwZJxU+CaZXd8BBfW1hCk
R0jwA0QHM9svjcY1ewsk7plJhnncmA00yaoDBNRh3ta12qAvKRe47nViB2RGyVAu6XJjcXB07GHI
SoDhA0JaE1w3+sAkyRuyMP5HOPC33NgGy+H322cAK366qCK4CTAsISalwlqqjcdkCLG9F51GT1z4
pp2ZEwsc+J8doxnU7pAPNrVrF0sZM5zWRHiuZVuwZkNtb6bcPKnyJXIQrF86M3ZrptR65hJcLq6b
rdEaNPjt7ibrTMulv5Q1CDDHa3/1QaR5lSC3Kgapvhnfj/SAjh8NmfqlTiyVvdJ5xZo3NnnJVJ3j
5qcOk8hsRmTlEXT24n/Gh1b/jz5tkA+PG6vS1n45EPLJK3rCRU8wGvS/km6dk5nmq65LyNLJtghr
is7B+KjwqdgW4E8Tsl6x+ycSrWkyT+cufKrR+/3YjPyd41u2+n51aSAo5blz28vluuMo8p7YSfzy
bIAwldNa/05jnPg7qqeCYLrSfLmVUckoLtdNXjsqPPbqNh9zNEUk01GaYg1AYKMJupmiPVGjMTLG
ubHi64pyvspDqC+sRrRpJNReqpVdpo1eZrjTPAxMSoiIMbGixPM5uHtaHAhl2VkYtm+AL4P9Gf7M
qQT6KoQjLYCWUZWj/F/fKZMNBJVPO/u3u4umn7uSLMeT2DGJbqQv9TZ42nSlvsoffXO04mXd5nZJ
/ama6KoKHlEKQES6n8bQfB+qNRaJjxT6eEIaJdYK4ucX1n2GGcSAsYLTWsfMcM+bxV7rYSVqrXEs
gbEanW7PUXwi2FAhYRDQQ33N9GqM9EnlYUadKzvrqoXUAp3Y+6xxyn+1h9y3ggfKKo/VaHTAwLYE
EfjQxHMJDSoaH9+yRUuWUHDMKR8FfpPrwALPT77zPGkbER/VQWTKsoOrGHkUme/U6MlHAC0L9jDV
vvY7BiSG9MlIj1u/dJIlMily8THEkrIwvsksWIUmUbMfnbAIJeVmq49lNUjAun8ukUWwaNE+cmxT
2Z9De4u7kzAV8E4Yyth8LATkB1Cwzx5rcXwJCo1e2lO/CcUKFgdqjm6qwvo+vOKYVAB4UnqaIHX7
Gp+6GZM/Jk9w5ME6PXANzi8B/NJZhoBS33lbHa5JtXDefznXOiqVymnFA+VDh6hDkmXQfwrgvYSn
nfWAf4qD81xOmKnpplg1AheZ263hB2isTB9P2hVbPzdK9N/IGI/dPf67onxd7M35J0qQnw6Pjf42
79asLS+qZcLq93qwJTJhziWWDYc/evCRMFsSsTvo3/VLM1GC0RlTDivNGWcSDpUPYneJMTeeDJI4
PxjLYb4zBStFfHjL1EoHX0gShqiMgC4hUJe/f7CrrSe/za7ywfLGvYtLGH5yQoy3zUGhAS+zQrCj
HYRdwBHl8vR+KC710ius4LoZw2hQ3TqHSC9JZnqNXje78fnDtFgRxcKRdhB/fzmbvqGp64o4F+Ff
VnC6GFWx4J7sN1LbfTKtsolITAK/lQr42q/K3ZQpHomSImbV1Yl/wE1dSiac//w3IrX0UwcTdSd8
93dvBDGQVqkrzm3Vt4iESFrhSWG3WhCM19AeMEPxrsCs7m5kAEyP22CZ1AqTOu4VaYJVuGZdqr3k
Pe3pwTz6qOlTlXB163FZMu2Yt5i3+RCaQm7LyWg6XcJQXultBc7m5OX7YWrSaiNpIZZeZvLJnmsE
D+2rAkujYbwYzDetvw6MIE5aDz7MCDO3tJnnjUUg/EkRCXyU45yruq8qPVNQNf41YhwMasB83mXk
E3pYNgOZPgccF/LkalhYXDVr6RhoW5UfhNk3v6IXjZjxM+PnMWse828qdLvKulpFej+MIsNh4Ou3
Gfoh5jisFHc+HID+QuXUsKUAp7MYL2tvJ7/HLvuemx9XpLYONvlXtK2UsfYq0bsY3CdKJnewpejA
493rXfKM0wS71EZNAENUmFkY/EaGlE2JA6ibs9Exg8hu1GofYXiWEqcRSyvPs6QEIlzOvSsbMd+K
LZbClRLrXKGs7PMDUqKgksQsJA00bYiSi5R4ZLMg/BQwFbQm78qVF9FsKNfqg/cplT4Of0h8LHqf
lxfBhRs0htqRvMRK0Nbzt5G/2jl/fBsu0bs6sjhxff3mogmC4iipIN5zvQ1p7pUDflQGvxr01yKz
zKbIeoLSt9BdTwOzXgoFv1abk9poy0UQoak5QgRM6ta91J6WmBU3uocLyQVfHk33RTL0aBkm/ges
RFIzk9pvoYm1wAtsArzjQFhpqPOf2wMWc+dU8ICOezddIK5v/QD4y6mh6AHBmv1dslKua6yLR6CE
+OC42dzbTmA0+JdqvumISjaeQ5bkUl3HydyBS8P10lf2VAyD91PJF3/WzGbrVh0laq/55eS9sm6k
lHbILgaOJFXbEXD4SIePeaypMv6LlU6LNPw8M+OV+qb6P2tDa/ykUYoX58c15pOLkgGTB4r2iYoR
ZH4HF1EImI/C6TUSRe0wfOgF2ytHjN+ymojGLKbA+IB1qRtqvc0nahrOlz5wHWVdTPgKJncsSBpN
BP4SKAe0uZVf6R+AS4MGvCPfMXgvveAMk1EqcfhGRSmQ3sPpbyZHWCNiSe9M7gfjAxcrRsxmjIZ1
R1XxrDoi/LG9bLuVHIG33xP1YYagUSsget4Kng6WIcKVJ+wgclHMfPYh3iH2EJablmXCdstyzmB+
pG3HW0r9PsrqLeVk/XVq80qP77uBT3/zpDWZW3/wcLVI2VkrG+p7A1Qzv1erPCdxcbjBHHsElGk6
FDWdIOwIlTs40ZFObnAuubVT7qUrBtWfXxiTkvWSulpz4g5HwqqD2xP84u8FpHYPRp1owezXpYpH
Kf64yf7khat7M1M4lL1AQjKtUuaRrhNpB0ncLvTFRfJveiv9lGCbqqkn4UUNkctkYnCOV+NXtzWk
QY5PZY/+Zi4J6andqKBZlOHTMsjs4juRRyOBX3BBXv4MRQgBcxW7KzWtPmu/KRIpHVpjWurl/59p
SPGnjGZNodxM+0/b7PMikEPb8EXRZDxcp5mBUDvaqdLAN/DchNQdbMOJdn9JWPr6Dm4nkrOKyWe1
Pv05D4fjgFc9RNrEvzhiOC5rr9ywNa6rj/YggodZ0U2lP+QG/EapbTiRCA5adSW8Y2QUtlbcG0tn
FozrrbQPOHeoMMb3l6BeGQyBruV6Z4lZCrGoIQDwi0xEY0RM1sw3tLMQom9krfHECb7Ln1OENHD4
AnmR/FQdcRNyC8LkyQrq8pqMfN9bQwn5jejFAVYtlKlRI3elBctzoG80LcORygc85SZDVHQZAmgf
llmG3PDxdX09IbbNGSvVKh5N4Mmwiz8S8FCzDs4Iz4qArDRdk46Gq59LOC95vWADg2RGDCfgxx17
tISqCEEwhK9ZcbEnRDBCqFoavGA/eNg7oAnAqqOIWjvD64o5uByB0VN2ikQiD05ezuaVKGPLZer+
WwXukluKi473IrT/qz/6uXNyQrTfdQQ65J5uJhjLDU5210UckyhIctHi4f2fmZfDi39UEuHTSS5B
f7siGqKnQI3E3/wnNiwiK9NjxPFP37RB2rbau2dck0xB9BN2lnkQR+jNR0knaDe1Uv9vZxiYQdlo
XtMLBW38PCfSPKGmVn9rlNKCskPUMHkEnj4uJwCTQ30Sh3mYcodoD63JgU9D1fd7z0L3tDUBGZXB
GCsOz2MqcEMhIoAcefYM+WplNJqHBH0ybOQK2UlZhJWmDK/c+76FpL5PABBGmLP9jwjCDXucocG+
jU+WT8BSfveYG61SHX+D3a1WamxhhzdYQcyFpf4fnhkKn5KPrk1DPhp7sjeIxQ4Ux955u5f9R6lX
d/g8kJaBCCcI2DRYLUgIC4z3koDYFl8G1SI95flOh33/j8OI7Nf37RrNHfg7zjFwhQA8RJQIX6wY
hjpCLs2ZO/KudBCdZKzYCwi1+v08RGSlCiLELATq+FOi6ky6el2hLJnTyka6Khhipq7TKoQxC8HW
0PIz2/iF4Vb/jhGF80UOIzQ5duJL+GLGoNI3jL/OpnZ7rGWF54kNg6z/CII+PHhRHjxJBiicETO6
ky/ClltgM5rmR0V6Y+5yfHw2VTKEiMSBxxagOgHkBViLrQDwIjsv+13mCRQMaEtOljyNVQr/cSCR
jzn4h9MZqIVlJbTSY38lfUz28wSTuylSjsHNb1lJ7WDMkdI9yzpjgeJ6XqtV+FSfZwKHgFP7+9KB
fxvmau26fQ0tcuT4EOJKQlkFcJs+iECOeZOhDm/OZIOdDyH4fO0AMYOiCg2DoN7taIXA67yuv46R
SEgTN2S2vxkDhEy8ev0v13i+J1WxeiW/+AL8VjN35NgTcAGCcTMhnTQOnZpieBfM7AeQ42cmSZtu
9iGrg7P8xaINFFyTtZ84vFjjiOGaM5pr80DlZCMxQCKxNGafnH11vMSSFZwVKWG6PWVeJaFjZOuw
Xw4eiXvFspyjSsP4hJOlyZCe96pnjVunApbHDqMO3Emn4Ib+5ID+Xkeib6ma32GwWtyCTurg5Wuf
6eVQR+jrxAr7GO4e0xg+9avSWdIFXodTJcx1KUwdETaDc1INRO5I8Td/dzDAC7SUSweby+BLequz
+RqsWVhRRwsdnWL1k6ti3iMUtINCjDG2onnrYzVT82CtZVP0LbkGRPDn3dnsmX7Nmv2yKTtmACPj
Seh9hW2K60hgTZS1+i4IR68eU9X/O91Jz3XD2ipr/j38/ytlM6FzVWda/6Hq8WF32+IzXGv6xcV7
jwtebH7Qr1Mm+cbV9znDMTiv68LUwZTTRbMb6bsliF0JFIonif+enp4/xiqxIWJohEhIEpFMsKY1
LiD1SjryW4jCwmYlcmsryYBbjr2t6dUbfYbX0StK5RZw8KjZmwF8LaZVt1JrGpO3qulxjbs55IJ/
NL83/uc7zMz4IuOJ+Owuzu48KJZveB//1ubANBNArjy32nveKeNoJOzVdmwCWX+XFUOiW8daasJb
JVOuTr6ad2hIAQXuGg6MzyN4a0MgOkuNJi4Q/mk8Z/8XxraRyPD5TbfR99H6II6XknEvB96790X4
1Capl8gIQ82KbZmY8tQ6KNNQ62IEh5cSxo2tBiHaVbclWj7s1Xg5MzDzd44V5KG0Xf+57NdL3a/9
0LfUVxrsDx4pGpjSRYrKtCQANLoM1U9Xgvux9q+OnbkjKWv3z1AkLaHCiRXZMkdqRXz/PHy1rALR
hSxqWk14EPbepklqBmudBcg2XSnWUYLh6UsMGWXDTMPt1s1QpmVi/cuFqdFT+5GnjiHgsX6qnYdZ
hImqMSY/4V45dlYQzv6I2co0wtmZrZs/32mYyjS/l/1ppeLfWz+DW2M18cT+aDU4mD2QdwFksT6K
jWx/qGYZf5ZBY+avPcaOw1N+8encPALO/uphHsd9WhvCYAjvzVhM9XXfvwyiW7VkyoeA8DYZL5yM
HtRZZNht1xt++cLH2rusTnaRcXMUwnOlIr71+uSlVmeii8E57ov2f2nJv+ubg7P7fLIOvSfdmFBU
3FcG+NvjUOUckc3oN+7RH6IwMwloBb+Yz4tg9C8MHgzlzYjfvk83bBbJszLuLc5EmQnCWcT+YYvl
CTl+gINj3on+hN72ZDix1xjumRijYMabdYkXS0W0xEqIjhsxN4akR3SVVtNpxEm7iLQUi7O4658o
PbixaOfyQvwHSF3cXm1kCjrZ89w6FE4lEPpEsOysr1rO78YTUNeMDsud2W7zEANskUmsb46cCeAN
9pJOvkKZwrbyPqGSkvsMIHXy7EAe4yl+HCEhQJ32t7ypNCNA+mUM3uQCqUD2WZhqmGUbn//TorIm
tUidYwlxRlus7/T4XbLwhxxuuolT9Huk4xkxpNt8/7Fcoa1gRwJ/7N9WApQIkj6l/vbbnwlIRWxK
2kiPzfUPA4cHwX67bPwt44LN5HSCJOgq+nmgfrDquelgHo/yti0QVNHi/eCQg9IUy0ZKAQv0pNFP
6hzDR05BWU/iUN0H1GPjwOb+YWMIhLczxkAB/u9noAgcfyFLGtCVBX0F9Mt5DnLiYiDBZCMlnByz
+fYts5kGzFCHkcciFwrueP/0W9X4PvdHjVorR7iDo8LCcUgHl4VYDyJVQC7T0jIqfwp7c/Rv2ppN
+cA3550hPoYypXhlWonun3yUkzRDVdhrxuDfsYPxQo8GjOPXgjjPuXvifrjZ/5XRvSHWNRfm2cJa
WBiNzz9BL7noSI+NR8vZDSemySJdfce4QIfdWHab05ydRdaI3/EIzLmZOMz/YKK19+3dTgR7N5tC
BosK7rN2dlU2mDAQd5WZKlQ5e0oGf0TkjY0iT/jzc+dFBfqScWxIFJ+y3fjHWWxMRLCV/IeXSVIY
csPNUCjx/CLEiba+1wQOsj6ZTbafaghf6nmlvLhfiCd/Im4h+J4HKi7hVJk4XosdoAaj7Mirm9Ty
4+fZieZaARvJvzNPiYOyOmeH4pdLdx8VIA3zr2i3aYsh4f5ZulVbqskoEGruhGpD4bw7tZ5vkNJ7
hHu5lNugkNvcArOxgycnFQghSRrvVNU+y+P9bDWJ5oFy0O7j4mEXdKuyRAD1yOnWmIxvt7bGokbt
3IyCYjuxKJ0aTiPNDJq9buOJV4/U5XTtrEF1X9tPbKpxJsebi7adCVwyC6WjVlkgckHeQGyLVKI0
XA3N/YQGGIkKbpdnosrjg4nld4ydwPJBaC9KaYWwQ5Y1BnXPlP3eDMUhumq9YpNn31GD3QuTFvH1
Ws3OHE3oR2cclV9uHgQjGaTPnL+sBnMmJQac4Ntg12cJAMZ2Hj5wdPCo4UEa8T25cRyRDuNnuZ9V
XTCN7eSWn9jV0/XFXzUj8Ssuro2uKK8D3ysnLYN5S8cyhSo5DLQxTy/UiRCjLgmqT+XJPhz56/91
8DSOyi/KD8v0CtNJChQR8ysUROmRcz6AFeplrmiNgRDaDZ31mvKigEI99MGP1roczVuhTcL64R8z
SJI5ull6pyN1pjsy35P/DJY8K2sfLiIrSo+fcyg26eQMTg5C7Tv8U17rfn5+YSc5JnOsJ8F/Pcdw
oTfS7xRtXL3AdufnRhvxGs8ISjPP7KdkoydGefxSdLiWqynNmQ7dtIXnMVLSFtC4RljysRngNa3/
Dnj8DJvgPhrjr8Yqf2iaFrcA7qOjU9fjGd1DKprk9QYfqDRQfaCME4GlK8DUY+85E1jy05db3ChD
vLscjgolJCcu8/d+t9r8+xBuvhkGjD5Zl3+QAwsGR4cnKpyzp4k7rpJIu1eLpnGvsfUvY1PgBHD2
VZMP5i6b+QO4kwEKornQkEGN9zp6eGeNNjeqm4oGHvQy4Tlc8PWjHUywNwfwZclKrznXiOT5e8fy
z/aLNQnSlob03cbwb1dmlb1HVkxcaLhVbkBFCOuSWSKl28jPZxBjtZIvGIEHs0hpEiR9ZrXCJ5AX
d6LUp0L6v+X33yv7csKnycvU8H+vRFXBIZV9JybT7AIo+skmT0DsvRidv1uf4v99h71h89Xe2w+x
OriaOcvexUA+y2o8G5yePjAXGt3kOgBxlRk/zZbfYSS9N74bB3tb4G71tiUN/As3N7jKFY19YAZX
WGfMuvSBkxrais0VpQ9dh/7bgfLuLk41fJXrUBN6dIFhL/13g9wYoGpoghfD6dX4NTMv8uA9jvQc
Wa4zl0oAOo20sqghpnYqR/HK4aXSTzBpL7BItVIqyqQ7jYgBqDuFtRO12PhUIzT8iLcdqlhcL38L
0IFGsxOLZDQQ2qmjtFDhFVziIXEFKch7/DKEitIrUW/pBkH+L6OzAD1VDo5b8MhW7+mxYQXGIAen
zkwVLySi+Cm13+T/fGKAdMrvX3q7Nzq23bQsdg+oLeWRlQN1PhbdeRzAs7K7I5KrJolO4r2txCRs
aq14sBNOn7zejNr3kWN74/JpjDjLqVwMaTsFyjqUbd5zTIG2zsRGDIiYXfao7zLBi+KXKx/Ao28q
fnoBiFkSUvyqlrKf8PainklXO+ayF/bhgbL0Gam5M3Yt1QY2HYYKw7KZML9MlEHfJgO2lOwuKl3B
RdwrdkhqAqeqVWUMwf4mPKGrgRACyRK3rQhmyOZh8MpSYgsfrVnighw20VtD2mcOhRunXhdmuJll
G+znDKviCYn40hOb1t5bX3o7dhwjC5JlKEPn08niB6AzdM/M0l+Rt1/zo1cXz8s9gH3hM3EB84eA
aP+StH2F/ACsCP9z9jbTv8gicPIRv8IpLcqzHCJOPGiwqU7PVL+fe5XLdKnDPpHFEizMhQ7vzK0H
RooLTcFdcZ0sZWP+sZYX7do6ziQADcHKmxlRz0WR+SW+vD9J0RpYjBAi03JLr3ONW1CMgPfB8Gro
3du/IxBasyQS71jcEkMsvhRvYu6aTFSK/IQFSwqsZc3pB/m2nOGDF0SExlxX+e5TDXbPt6vdIu5Y
XzQSzngXuy6RAdV+aBYUloi00qVJciMGur64+OyzxP7ceAyYPcMV955irWDs2fX12dXoSpfCH/qs
6QDZ8onzhPch70Wk4xYfbBxWA7deWxJlQHGgb3LgOv2nDMW22lm8rVzd1jbtpkVG3vCSC0C+mwOw
kHlLn5D0cu6g+xErv9U3UC5KxN1Od9Tj7M3fkh99KhrrUCxMjx+HevmOnjUrbcvcUVjbwd/IkvYE
aNo1sS7OlcpLgcCcFMjzMRPRSYUdvXFzQYXIdETuLYG5GXTy2Pt+oWOJhV4KN3M22ZAIilpoQlSQ
xgtNS8t2m84uPIyJzf3G4eFti37ctmyzzXPzLNg5ZvmT1t5LDGTOZzQzPxylsKR5ixmI78SCsaK4
9PczIXiCCswaNYffbQfDCiOR9T4PQvkeunlV3Xl/v+lG79arDZ8N8RwZufxOnaOR2EzUoJEWD3Xw
3ZnxDzkmqodJArZoHeqYD1qMxBGCX6SWMwoIyqx8RLX0VtObLA3pTA5nRrLFsxQm9Kc4P1NiRAOW
iW6xpGlMGupgyi4SvVGgVBzTg1FENbGDMHNOq93lJaVgv8oEdslzcLxT5cFibVhWPC90wjueqcC5
IsF5Bk0mU75Q03KgB9J3/i7X7cWeNGg27Usb2ZXpyLLpMHEyW06Wi6A+Ilog5mjmK9UJm6II5zWv
I/2yPP1RjU72BzRuz54GnVaSg7ImjxOyA+2/46TncbRyCAkO0I/g6/tAjoguezzjFeXmBVM/TuxU
ex6qlsnEE6zahNq5lUJhndUm6/1rWyxY7cX2XgLWvz8hMyVIEXtHfbf+S94CgUifZrYK6xHNjblr
emCjjgoAXzGtkA4EE/YwJKsGNKffYxdBr4t3cQdkMd/4GQw8ut+33JJK5nfyoiwJsZmluiHRJbpx
U1DHAm2cr5/6eTXiX6pSMUqvyhb5Pyujf37PQXpj93UN1CrvZLbESvZJbyN8Ff+zHz+JrFZGiBqs
8gc7KJt7wDZ54ZIzJDlAhwcD1iq5Pv54K6NiV1X16aEGCjyeEwHBRImRgxvEtn9bS8rzQQQfs5Eo
bOyOIL2EIN/OCt/F/y4WnV1g4m5RLJBh0b4afQ0TXEvO5sz/vv3S8NjEmq1NV3QbtP5rTl0nFJRa
CNafn2wkLUhcpzG2XMe1+m61gl8MvfEgJ2Hep8RBa7P9x8v3/gn+b1T7FXsgukMNAQM70QLFGnO/
GYH/m4YtD2kI1b35IoCGXCi0Zcpq9R2PPE0q+SzFuLBI9dKQXkDTD+JVRu0Y2+yAgWbqgSRzD9Ze
GqI5yW0qYixfJfSOklUbLmE0ze33Ic6YnhTIDPyXABGE9QDV1ppPilKmENspEg5vH/hcqNvBKf2I
mpUapViYI5b0c84v/MoebpBsgzIShiR6KUo36bZBhpMlJKiwOB8R05Vylp3G6+DeaM/q80yevK78
IXCNG0dCg2tpDbcWK0WknfCdxu883zjgJmCEagBsereceJr1JBlCfxll4PwvtNMx+BY7Q2T3c99R
K0k+pESBKC/6MpgTCUSElyvV3Psr/Iiw/8BmZR3mY9Q4fe9uI5ajn4+mPjzncZAc/VOXpaP85Vwi
CfN8KRH/ZkoM+XcluM2JaoAviUrTxXNYSwXX2QQoXqRcBoQh7VhE+Jjf+7H1GMUYQ78ypkmE0/EB
1VGzt3QIfIyt/aDhfyIXb12E6Z0CLV76cO4ar0j2KSOeKtgJfL1ZIb78xDk5JyG8ierkHHTn9k2w
qVd8FDX/SzDeNFtekEmDXplwMrOfyQDw6aUbBVyvuDXM47t6FqyQKP0ZUjyn7z+oVrCLIPdiJ6Zw
HzWx7MBcXSQ0N4aqsB7/Q9JtZ1YTC6GKH8bzH8hgBvGiWFsaH5uG+Ge+DC5GhxjzwPkMLRxF8Pu9
0TDRvflNF/l68QyEnis/TS1f4K8qMRff+kQn3ClWCNtGrSWJPh0R5MsjdG+FRowOQk6hugV2dmdg
sIr+7aLYNq7B5qEZjMYZsXtPKfjiYQIC7YAE6unymBD++qL4ML6zqY25inZZFU0Mr2uVdyDX5Ta2
OCn42if3yqylWGVrTf1VSNT2sJqsFQa38zRkSooYOeYeNSAfWvcJ1uDyTb8LXm+o62jDea7AJXus
sP8AFOHFptVp8+hxi0/KLMw3ziEaPjjVQ9R90Vj6V4MS7noGbIlH+prwbswvH7f9Qea6ubEZ0Y75
MDDs4FbPAl1NvUb+P5s2/1iJpPThEKLbm3OH1mI6WRcGAkRagB9+Tn4rpFqJStQSiCqaDbwAcnTb
fDptjAvXXMsdzbDz/y/KeaG4BelThprMJ7xUPWf2RJoz2kdIkl/KsfRXt6RE3gIjqC15nhb4DuqG
SN2GOb9Gs6ParwIjjsOZiq7GMsxtkilll4SstBZqoUD6WXsgDCgmas8wPQwqAAU+AZHUPJRvKzxi
EG8avbknpGFObTZFXPHOJKafMXtkYgFtJWsMq82dvbC/4ipM3P9yLqvhN8QtGD4PyO/YKmdF4ZJQ
U2YHfCV25G1sgzOatqm0hcj5Db7q/cvh+RFLqQR91nou1lGt29Ui+RmJJ9sLJNJ13e2Cag3tSMnf
uOz/QHh8vleC1HnXtKFFR1WiBoF8FMmuOEoo9tlhs5OEi5crATgCopwRxeuWplGOLErNRz8krilE
3yOy5wBp8x/WN1skf2SliZtc7FAUk874VoBrz9hDxRS2Udpx0YHeFNbqoPvlTSTxvOsLChW/ZE4Z
fSsJriPSBfpYFTajfXheo+lA5jsnX7TcD2XKSfFPKGs0y/HL+QmwQwsPENhUW7bA6AzdQKqSlEAj
ytcnzMt0rOucN3NwI/3fg5BFcmStIvtAtKSynH/60rkXx8dG4GZ2WWiRrk3yb+EYXuP8jcyokKu8
w6CgHFbj/1zv7DZSficDmlZFnkdb1EN18/gjd094RgYGhlJtxNCBd5TWgjWUEBGvyrfCpvLw6DLU
4lepzJAnvvkUAafhzBTjEZNI8f62/OKcuGhKomisy8n26JOf/p/FbiXhtKPVgZMnv1i4tn7SztXO
NsGvuYXlow1IzWCXmQHWfeeRrcakmx3gK/0SQYBoE2u38s4115ZM3TAzqBYR7NHmAk+FnMFYjQ9A
Cpn4NKItsbR9g59shGR/XFRXaU1Q8rCK+abe6McsCvdaUdjb+sZeDxqdhEzG2yTyw1vGIWSA+OPf
pgASlbAVJX7dhyySZbvT6M9JD8TZFm0ZZfW7LLJgqTc/uxxnoXBKcG59jI7YgXukx9SJBLwkLtbA
1VMv4sgN0U/1lBxbayz6iBcfgdo9X5A6BYoh6YQ1AIbl9dSuqIfY9nryVmqbU1iW3KSV+OQl4/TR
e1VW5tRRJms36VXMeNievubvcTRQSnKj7NnlvXOJziqkOeK3EM/rl3GuTxHMNCAO762HN+oUJ34l
bytYQItBeOzmcAKltKrLhK6da8OLwo1bvq9e4Fp1PSnWWzIQ+Uv3fcLfTywmYHmk0oiZ7JHYmegR
6BzcH8BcuqD/NRAsE9Hhbw8+bY1Ee3lapR73fy2vDJdmBJ3RRJHu2z7uVpNK5WC3iUwntnIm+6hX
1dMdILEKJ28seG4ss89gCH9UI/Mgdj6xoybNLcjo7sg/ouibgOKcrUlQjScjmUg//xMYNzmCUCQH
QqFFpYvu/7VJAEe6soDyStW/duBSlPLVLq0KleO6bx2eiHBY/P/phWu7hBIrS/CVKpkHM+hy9+Qf
RvmM4C4+3z0Godk3USqLx7M3NTwe4Nu5FT4+39lt0Q4KZIZxn5WnjymeZvaQcN6ObESUUtQ/pNBN
jSPmSFFdJtr1eWy8JSovg4702uIRXq9atFb9IzRfB+CJfOrE1FN0hYXMV4chBni3+e0Rs7tdLOQ2
T4Oy3hB8mq7IocCRQVBeHcMX0OiEFEVLLC+Oi4MD4sriIwrZJtiaCz5ZNErqmmkS8uS2pjCuXQDs
QcURipx7KxtMg5TBIdv+6jnIphNGBah7UCp2M9/4uxUB24CSRgwgeDFpdCl45lmmgalm/xDgotwn
rSBLLJTXBGNxMpsfDwwO8zhRnR4IAZb8sYC8mpQjdpXAixjURNZowN7UkNcjopPc/LpVO51Kkuc0
No07cw1ERiwCGNT0PC9D7oGJKnEcE/dlNn0x6AvChVAwAPHpIfdG2U7O7fOPivSI+1z1YOWDDR2S
9E/cPlc1sZPYp+J1rpJ+SfSil3di3D2lNhEvxGhmR7WL/gStM30vFmyEXvj2X6WtzaV2IhJpRkXD
Kdaj3UjxAmnXP9h0HtVznuPvtGKW16+7/wilSk+s3UUQi0n62eYLH/Blo6wCUG0n6SkmriSMgUjk
kYjeTizACTUcWILlDRRJUXxf/I9ut4x6DTzNQ/WDWEl+G5Z6tjqM6e0RbL4G0vkRNLYkR7Vz45Oy
9A0pQnsyHlY7NvMeQEiybFrsFQCzrB2vad2MAd3oo7EEnvAbXrrLNyySWb4fLsmhRJ/IXoEe6nbk
pom5SqgKLT9h4/1CpsgktnYnsemfvNr/rqIqlWZ9CjoAoePLluJXmlGFMX71iJdPwiYp+TjCNndZ
2R3YHLboUCVCFVAbJIeoZwd5pNWVcP2Wi+YKSgNG3AwhEc4tnyq5FbAomnWidDRFvE0ouZwtKH4e
VHYCzw+6IGGdqThnxzwmAO/+K5daoXlVx4uKeuN+nauyQLUOK/X3NSINdb97+HsM4bvwOqy3FhuC
vrO1laCRYwJ+0nsoXKMxi6eIGDkTuzt7MpQX9fVq9xtAN7d9bRWlQ8EREKpLQ3kMYLDqHoyUKNUl
xVnLmZzWYasPGRbMLmPvPN5sq2iOolHrJ0M6JFidL285gHfSIpMN/7Ry9DzWVmPc7y74tGnEVqZF
CCTjE3VtvGyPgB+UUxXF0lD0Sm6MwppNwljgrIHTlOxDC8b2xfog50tsoUm5TlHfvQTYIpLKqH4V
rR4lGas8s/cqN/FVmXgLLhc7sZKsM7PsWSkls1OaFCrhy4ZykPe+AKxQq9tyJDd8w1L7j+IHNvut
5DaTmmbGn7jKa52FiVd6iMDkNM5Vp3hFF7O5+/wRBeOMgp79o842l2oJKlUfrOBNV4AuqiX/Wi+B
GQ1U3QR3BooAV7fR0Yp0n5T7ALMY+cbihC4cuum2dV1z5Ipxa4aTP6KgNW1HnBh8eFqh6iYbOBxI
Ho/FNQasD19FWFSRD6xKaMIm9v/jyS7HzBo6DCf58BUls/c/2G8DSI9JT9szivAap5bfsHHGgWsG
tRvGAzR581mHhaqKjSGX+1AFK1CH2ddBYpS6WcTvYdi/SimNratz8sWf1AmBOF4R624+iOUkAdPn
TKtZXBjekAYNVv//1RPJx2URSTSp9aTPzD578TcLmbe/IfgiD7qgBuFqJlVVeQtsEGpLgbiCgGNX
3i7k5i+tMZ55IiaWDg6eWRK2zN8xNJjSiSCQ1sGrKdM/lSHGChkHYgnmtTmFHgjWlxXYFPoWUQCf
rpEuCvZ28ZvxaC7Z5YOo27BZti+T+Np0SF2+pKRbZvUOgab0r3HAcHgRm22dVFuozel1mWPsZsJ3
tiZwHCMZ5LE+wh3jpEhHIFjs99Nk03OlBmfH/5PdnkbKbu/vU9FA3SU/TpWSpEoQ+IBSeWBfSJBc
hn7hjxGf1dcyVrzK3x+FnGymAgW4kOABUUQfe5KwKC2FSD59j6TxzD1pqry7EkA/u2yai3NwQXPW
tYA+hrIw3w0qxr+jr5OgTl61WVW+o4mn1BzKnJYyH85D/qr5Bn9FzkaBK79lhy8RmofJ4TU1fvHP
Ka+9jq6FOKsT+Ezxh757AUngX8ZdXB3c0wGTzjgGogg3hiAGYHJzz3MuNSiq8yv5kFX1PvCJIc6z
N0sjcIsP5hdE74LjpggtTD+V+Tug6/f6qIE5oEY4yt9lBTxYS90DBV5dsvu51hOTltSbY+kjElT1
/9TT9c3uH9S4UVctj7g5PG9WLIJw3QmoL/kHlAQdfhZQFkypjlv3WqN9d1wfdI0rKf7yXoOus2Oc
YGRiaFfVrP1S/vnSDYNX8eWTqAqPsC5AGQAxwR9whKMYIEg/3sr8ppoMmvSvVACEVp7DRpEavyJw
qA+n8jS7eZx5rzrd3otctbPYT3/gL6Y/QW9W4DO5th2oJlClMVTrosfmG63AIWea7vKprt+d7stu
7DMQlHn2uj7G6z4RMe02YYPcY8kERtT6S3VwLYz/WVvvXFUSw7w3B5ombvKMYQal7Rn05WseWSYk
45ASiUnrVy0wpnhjYxGViFc8StZpRkYdfmbooGoCQrULMnh6SHiW+DyIJxczJuHRwFHH39hs+ZH0
5RByi65RXXQ9F9/ZyfWX5B8F9UFQ2Q4+4SKESrGrRbxDkZuQvJ3LYnEEicrF/TppsdcR22myubaw
ddVQt2oDh8ptUS99jj6w0VPnfIVLWT7bkjw6nqsoF6P1rm/s+0+Yqm9Rv81RtC6pfI/HMzqpdGvH
D9NbtgbIKPnzZBwIQ91gm7od/E23K2J8xpSRTN8fgAmTwu89K2732z28HM6i2QbAMAj9wTtfNypT
cNAZcN9poQNGcgTR/oo81QQOvn+OTs+SYCUhnHInDYzQRLC2EISONb2okDxvlzkzP3OzQE/iFGjc
jeHuS3klUxtD5fqYDWuaCjfV+GvkwaEublKFravFSZkuVHed/cZvAi7Lb1te3OeuqT1Q9BwoUSKx
QGFVEh0J2un3o9MD1k/XT1CbsrDSWkSWwevLN1nbBxaKkQDmYuaNi1UMBAIH/ChDoGboQVs0deQg
mESiAIPEBvaR6vgBvjPEIN0qIcabZb+WIU7mtfB8Aq+JrJC+4XWFAKrIzDchFQDqxi1qGBOKXl3R
ByVVeykUoP9C5e2Q4CWOUeiSa97ZhtFweJXrYQqtuNj+jzvtdIZKkx4DOlPLg2ENOBBlskUf1Gfd
iTsz7pZ+GcSXLBPorCVbY/Ruzoa4pfvQWd7micRWih58UiXLEmN1pd5fAHgehD3Zpib4okm/mGGe
0RojHwr84JAKHSF7nc/UbqF5Hg6MaidpjvbmqXsin58W5K4smwBkt87/VT6SYuW7pqSQun/QarA0
cFNEU1gtqoUGKuJcXHI/jVOsVxI1mj36VAPrKYUwACExgV1FYXanSscu3dzxHDJD4nu23980FK5e
FMXvKkVYZI7eMe5z//vj3F4VwCPgDg3PAKQIiWoGkL1xv8SDfOztzJoEEFrdr5XwPj+8zyyXtGdU
gWLVRQXPvgSMc9s/VcY2PGVwRjWS+rm+hcZj0pBBECN84r111cBa310hPOJpabEWradnWpb+uoFb
+mX3UUNucTEyAr3aU+9j5GOKNIhkHBTmvuYrPTVeVhSuXYIkXBGVZi/gbSKTsNrQ1TG3dScto7FQ
2w+PrwTSU9WYgNSERwxfFHtu3fx0PYj5wN03ch/8EkdyOqXQGPTO2nCBeusKlA9ueEnQ2Yf4Pzt+
6lg66y03HDrfTF4tClqEO+r8Opz/rHSqjaF/WGuqvLyl2MSnXj+Q0iub0lqG17zbPdDnMdoDvZvt
jt4fQiqcRKsRa2GASctvlUhcNyFWvfuDYdmBIRUNejnI/wcYePvdBKNU0egU+8RisoYVjg8ZDSXA
iHoOvsaeZsmVP35W/wz1kAksYgbcsC9yiVxqO2ArOQe5+v8E8dcslrwdr0kwGCKP2W92kyq68pDN
6mqm/ak73xdhYIV+TATemnpULrSpjhHg+aEgKLcdtYeETFJukwX5hSAzTN8Fdee20IO9hxIGJwkl
0TP56a7xzGQ//TdudYpYbHrRfKT+U+rvXol6oA+e7JKJ7BTrkuBASWjNcXA7dnLg2QA0aX1mNcRC
jloRe8f/n6oExdfcp+DxKGbKW5N6Toomd+wS3ovcM5korZrkynWZsQv73LjdiBxVQby854ZnT9FB
Hf2f/ZptLxrD79rb/RkhxDHtScvDmeYNH8zHh6iDoBJZ2AOufttt+x6IcDf4K1NQ0PnC16T4fz9S
7T1uhxZN1INuieCpzS6StnCVtgSg4XruGsO035g4lgDIiWLo4jOUy26Rakv/61EZ0wP8PGUKILC1
/lIZIexjhdtUfT2ItGsWx66peEj6xq0S/iep1dLkEmdTxUeZ+Fz09cdawhqoWmwP2/HM9sbrviDP
wbWMwtmzqoqDIWHstGZ2qBqAt+UKYGTPk2lu0f3E10yEvHeH2GlLc1yrFUQGiXXzbDSyfBEG5WWn
6FirEtyeD90avcwewMxCxr0rHURJdYM0vIOQqm8Ki/aKew1nmoKvnY+UB5vpbMenWMf91DsHoSKc
naQMQ7WmYt+yZ6x6QWyBlqlXlquZm8jFsvABmw7bAe37zpz6aEgmivNg73zg4grR6YY+bIXemTnE
7J33HelDiFwPGgoA69xV/9+tSDNLLhgUH6wzk5dbdmltRxmPbA516MdhTYm5D62ZbTyRzOsiiaU0
tNQi895rMzcHmtn/JPAiKBn4cHAdrY4Rpj3B6923FHNXlvip8Igqq9TNbbYiGME0MwLKLZ2eCkgs
xYg4k/cEsrSN7VDh5sQxrkH6UBmzbhekxRz3jbIHKI6EQxNEcFIleEDl0C53dlW1czyrwVehuYLb
hnTj2HbhlgQZNnV0Xq2Bu7vTwKOQVibdKVLfHKzIkb/F6X3iYoXYAavstOBZp+zo4G0dcbIa++b9
X9tOJyQPAPkfKFf8yDJelH4IWd061WiJLeogDrZrYhOyHTxC8uqRLzLTos+FTnBYRZy3QyrFGuuT
tqjR/5E2lKg6jU+lM1TArNhiMotKiUtyu6aJ4svPe9Cwq4BPRZ3SbS8A9ONggjfgkeRCKIoN+HPb
ykqvuRIzHOyKH99dxg6QcHv7Jjuyzm4tuPpE0s2532MAldz0c9R2QwOH4JxtE137m+dBMsWrH6LM
y3qXoCEYlrn2SU8/6jYty8eAaMm+1anilzFNMkufpqaHoPbe6+oMzTZYONBxJc8JdnC0bjaJdNZ2
MlSuFxzPFBZW7NTKFxtd3fCEh2LN0FXDiOyj92n3A6igJtjnqvp2AcA5F1//qfh1kYciArLkYH80
OaoPtDBCf2qZa41YgHTPMevg5a4X+XopoDpOQNmvvaQnknRXA653v8TSICUhAs0sdhNinqSTwhUY
zbJn9ZLYoxzoIHNIMlOHnSQYjvDphnlB+THLq2ujZ1VdbcSeg67vrZeWa9bxE7qiGUy2ZzSksz+b
Hs/N29qGAzlY8f4XknI2bU6i7oonLWBzCO6Bo+MjaIg4UyHcKlqLpnBU4lMFxut9qeSqwKFR8T0a
Zdh/ASoa7dF2d8W67ggTgGREOVjtyv7vr86dv0vIDuM5H6wycyndJJs1v5vBDt14ZedhQ321bsaf
xICk2RIrGQXPWLsGou5lEjdj47CycsI8qluk+a6iFX8GuZSkRP4quux6M8K7PSPR3uHDs0nWJ0Fd
FGhR/TM1AvihTFhmRvpu43Vcr+wv93ZhLUdCcUD6raMrKF5hDW8dw2YzY9t7TRQTQoXzN/5FX0jQ
/ZAyfYDY4FeFLeILXciOcpKSAMc1/WOHAdN3bmmNnr6ezFGHbyL2uyBi1GdJfB5KW8b2OFtwN0Go
UcqQmkC7Gq6Dv0MUrMO8sNWCHn7lJnapbZM6jjzMgYLrxQa2gyrKShPc+e/86X7aR6QJTA4N6N1g
Qg+Y/g3lAC6ZWJX7CUkoNHdkj7KoDSPV4W1al72bwTQ3CVmtcAQJ0ljuH433sgr8Swvy8xp8VrK7
ttj4G/OdLWf5yvKBhD3OwbQaqaDt8k6O9J4huWqNs4hQvvU+uN+MreQz/LC5mUE8zIkJNC6xqdqc
7r2DMnzzFmA0vSWUzP4n4OxgeWn8hTv3FPT8KQuTJ+60/Gma4cP+jz+rfODoVNP5LmBCIEX/z2Ez
OQdhWiV4jYDFjIzOemVXRu34lh8qM1w6UpcFVqJJBKKyjilhy0xl6nrF4fTC9liloK6kJRLpWkzS
x7kr5V3txZJezH6HBAtBW3k/3aAPtHcBFqMWrTc18rLYnXr2hiPNl6kqzNpBgGwvAV0PsNTM8+7S
Jne2uiGVQlFugTZrc/FrwHJbir7PY9Bfg6tRbdYJrQqm2sJNRSxNDdUCcuj0ujPpo9PQtb5mDK+K
TZW1iU6BbV0FffizQhmctnb8zBkaKrUsd+9QDn1+Q7HwR+9K21/1nmu0Ka4ObnTGCl7E3fYvBjdr
dPTcs1CXiKq5WiWKWBmmhSmxS81sqt9MXbPXDdsdG2qH+GLb8gBhCitDwfGySTdYyhlMEKSVwDps
RWtBImcUaOeQ/ehpsVaRK0VY8GMt3oMhGA5vjdPieoFxwalZm57F790T82/FV43vY+xSoXdpb1sk
a1OC/mKk76gWDyLpMUFpZlCemhgSMES5+qoAyIAjFvGGA2yG5YPA/l5YOROR6Y4+BQA0NdGMK73d
Cco5HuXEyhD2NsrGSY+s2WfoVNn42wGmhvWTL6TlhKpOf5qdX7NvTUtksxmVBwaAbri/TQcITrDv
Yd9sr6u73QsyXyudv4UyikOl5Qh7TKN0wLY3KJace7jBjZJ2fbVUl2EPimXXUvltlrhxwRuHDYkO
WtP2qeFp3do9VlOHjkGRpxtFzQK7JAm7YGJnBsegofFEUmzZBuReV/7SeqipWopFDP51dKQCmiO8
Bm3+Uh1ZgSfdv151X1xJjkr3RXEVqHz/2bgE3MhLhXK1Sn3dJ29Sf29SVSENjQ1H5k2HnPpEWNXt
YCQl6hYMu57NUoapHdgLuk0pi/GhI5Rxlndgi0FrvubMUWJXGF53yD1kOHWGAXqEipuxPvEQMY06
KCfe0dwh5u8iXAVplPRYRxoXM1//UUAvbXL2mYz8VzSEmULcqszsZjOsPkWfqVI1OjfeAd6f4RbV
pMTYv9u8zEXJh4D4Jyml1JXWFScRR1cLSAb8cVGDzCApqR7T6mkeprxyE3jfYTWvJ0p6hS6XUOtV
2cauGpYeD2q7T62PhkToThoN+Y0R5X+8R6gHVAD4Le7nHb/0WQoup3gzfiU/DO9BPW8VBo8eqnmX
QuLmC/QF9pvdOaSFZBFPj8s7RYMg5YzUCWOVZGaMp+vB5DcCV/aHmrcMyt5TrnMLKlIEIsIxK2ba
iXgpZrQVj1xHFaaKBYQ5ecFQUGGDIcVYJYpmRiqvwG8HSLNx6snK34aoVJfdCGSTVN49tGGyPc+1
GIq/6iBCdsl9ljECRs4fa35hUfHCeVn3BYnYAJ6I64gMC6h3N2BtLJqex7IVYfnpBZJSX1hJEwPk
UBRBTevloTSFU9ArHvjfBwGJeZQ0hW3Jg8ZzE0ra135HqLKzD8tjsTs8/dHZMNb9hMluuUg3otxy
kLu00J0guykHV4o5Y2z2jEbPv1j9KwS8y5I7YOMNr3F4JDVleFnsRp0PgrAnlUZk8eFlD9IkEMLY
zcIAE+KX77QGezgf7VmUBvpwFgEGIXJu2t4H94ohwS1o50ev9RPSyZomCYM6GkRQr1UdE86XVwrM
gFfET+Lqz0MKnnIL0vZzWk3myJf2peJx24Ft96J1lk+FGFPUZkwBwMOhabSpGJzs6vOQV0QB2GRv
khVaXqdDp8A14OkYF7IlidupwvMggvkaQClP3LORO29vfv21ie8KnWJTZ6tQlGggPZNsTazIYNaQ
iZoO0DZuva3BIW9kbso9q5I4PDeHIRcZAAaILIXS/VLlp6iBK/+zU7TEcw5lG/ZAh1AZo/UFzHPE
bPMPK1FjqCj+PLY2FGznMuBUWpe+pOCsUttqSrFuuF1uBjzhvRYyFxDqE9AA9lQ8cVyvyaSXkfmD
Zbm/gAhGydOzK3jqdPw26MEMJO7W2kaA5F3qU0r+8ouMYg3Aqm1iaIsoBw4VVhwvD/865wFAAKBk
kTxKUQsgprxTyY07VD2uyHKzavoSM9htXCa1XZW+0x3u4BSOTD8qMfo7eMLRUrD2LqJXmkikMgFS
fYNFeZJxKzeHz0xOrdLOEZ/FU47xncDUK9UZ3y+QBuBuMfHU1iRaaSm/fOqgN49dFIHqa3mXB6Lu
TFBscfRq0w1jkmBO5eIy2C9J2NoJFUK9t9NdrqywszqBDR08KLuVcMECL7OPuRUHSFSbi2QaFz9q
WdUFMeGV4IzuPfjUmYv9++mRCK0fp5rxQC5CAx9kTaJjeeKE/EE2/91IBKIHZ9nZAGT2/nwpeifl
jWHahU8b1mHYFF/5jClFkzTQnt8+yuGV1j267bXU/C8jrhOz/EgxcxAG/oaUIUH3fN5yn4D+Ycku
WbqBm8tUEFZtiKdJfKXob2C3fb8RSKcTFNiWsPlQk/GqrqIoXxphEqvxBQZw4FMcGx9BA603OwRh
UB2Ymlee3HeylDlT38guPzApt6RZuwThel3s6dgNMl8jUnAXXw0ZyjZeBvMpu5xbHkAJhQs33ZWC
BLXUb0PRAoSP4BrHhcuap4t1Nkz6SkezMP1CTH2PHwv3cOgW779z9de5KXwNvuENYavC0WUqTMxM
7H3qxWAcjQYG7SJ+hBQ6e2PXHl5adSDGCw7lqCfUI5+jVz1PHib0TS0hBJ14AdPEMTojNXGZT+PC
ri+y7wp2zosPCH9MmYR8NNyayEH9VXExrOsEFdQWVd+Cg3uiaOJd/u+z7pUeyN1Cb1hcLeiVSvL/
QwewU9hL8RWk9EwCprFvBc9FIAvgH8iucX9618w6KGAEIzli9vzYlMM1yzyqCdScrICq69JNd+s5
ImsoIIoHFVZdq4pASISqzIHdzwqazmmwFzWpj9Rct/S7oKTzSIngRDCVDEdsbuK11gAJoTJrUVYc
e/PhauC4XdxBFSO79AFmNmP2nBI1S6w3JsudnDrIuOqhEhYF0kRJ/o79b2PQK2Mv1bYgxw5K3bby
GSZAkoGJasCvemb4I3qERoD0X55blUbG0yHtHAvb0HNAcDEiAr99Z0F6yE9XiqjxZzshmVcJryft
fiWhEWhYgkTIYR5eXDzdE+a74thj85l7oQ8F10J6Jz8yGih7r1nr7nhQHgz8uTesjV7PWgMGjq99
SEpcBriq1SjP5COdQaFotG/OKG/DoGJ64bRYFyjvISUBxVb7hmlOTwQZF+59nUtBtnVMGoa3LHPG
BUEseAAaJwuQIxetVAj8I7PAS8PSFXWf5IrcpPSY86xfYp81utJXmv4NjxWt/dImp7ndxFneRcW1
hi0s3ghxha/7UPHbnfFsRCYX0Bj03dLBmiDBw2FlG523npvJ3WQkQUhUQx4PEow3TYRqf5e9uf5V
NuRdZNIlbYcJnm1MbU7f5PBmLSYwHRJ237Bip8iVFcBtFac2h9EiLY7bryLDouHXI/7LAkxLvCtS
jduzshRT5ugESPuPNam7dccrbh6tYENcjt8gPj8k5D4TahsByM7XtqtnegeOh/E3m7q8kLeJxUCs
5UYg0GO2sRbyobxwj2r9FkhcPJkhYkRkcPS3kTUW8bfn2aygKIjj75xZN3nKgpRdc7FCLnRI6Ban
OJh7K5ZQh81ofjZKNFv+6xNNOWLj5uSQn3JIsXsKSC7d/7xi6SSUDGe5geSGKaZiVtanYIAfCOGZ
B/Ddy/qIXXLpAA39oq7v0sHRtFew+MqYsHmxVyo+JQKWG+yEh6fAGDEYK24e30KkZSiuWo3LDrXt
PR5otR6fcxOBzeD0Y3+5Po7L+0EYOvtjpOKi02W3Jd5xsDCurIhCiWRkhR6dAziCpsf7yeD9kvV0
tfc77ULrhgOr7trIWcWIlyJbzzhg65qU2Xk/rKz33n1rY4wHUx1DzxYJzMwGfckd9DSVDyNiZLmq
Pd1dx1BI7T8Dqs3SO3grK33YtmTfJJVNo79vAd59zAxssVljzodQO5/677Qdx/UX3WMGi4uj8d8U
ojQipzbPY3GzrEbP4TVG2cGl34DBgpo9GPpQpmaRUhhaga2gl4ciq8ky1D81n+c8QSAmEIFzh8g3
Vk0tWKnVnlHTjFxIFubwdKoID6S9dStgPZEQRbvNxF4zZvNPwXeC86fZuoeYUMhjQ/VfgHnYQPwR
Rqk++vkvn8lYN+Gs783mQsaQcP4kt4Syj9/gK5pCsd7RCVKQdP/fCqfkTBzaPgqpLYoLYxKWANqg
Rh7Bzu2MjNn97Hab+ku4Ss5I9ZBUKBVJv3J6SwY3Kcb26V4kSQQdQi90hzuYJCDRWtHtD/W1u/uI
yV5itN9bG26caYRbVtWluQho8GU2XGLWQk8znEKJCTaMKHawzu8ED5yrgcEa6hF9HULbWK8Ew/NE
/dzEuZOoY2ZXzFed1D5aXqzqATfPTZxSz2hzwL5aEe5eCeRmz4OVyyzXra6a/5esbNlIFaF24LUF
DprZ9/1jf94wdJprYlmxpZA/JbV8c+zVZNNQqOu22CimaeqjjPCH4Alng9hkFUfmhhml6kR91V9V
hIMmtoKrcK+r+wRkCekqyiDZLnUFnwqhGSjy5MajUmwsIxmQau38etLo/TDEkpi96nSpOzn4MxZg
lLX7Lo7pQ+X/7kqjN3OuM7d/Szo++Zeo+mjwe+Vpe6PpkQ7Yb9uCcPf4wYtbrguJ9+V9O3ZDbefO
SdO/AHqLIA4ENZIQ+IUT81q4bNSixKutN3928B4N3yhjZJN1AYhbmi1TOiqr5k/0QSbdAo65XVi6
lrKxQVY62LkAUlWngjALHSBOwqo6lQikuq+vo8mkTBPWtCj115fQnTQ1vamo+mLo6qYUMTQi3swh
fccYOgCK0hzej7UGcJH/Avzniz154u2loaCJW+EdgmXWhtMXE4cL3zkXO0TlYgXWBfZSvzKL+vtc
NxqJYWdTTMNd40tb22ut9+leRhoWB2WLsY9pAmknnN9HmdRTj4NiJEH/11qGn1pAdK77h+sLieY8
Km0Caprfg5YKMcS/NiUH9woa8Zj491ZgTcrY2DYiZlISCvFXa+sCV+MlZbVsea8njQrwGGhzF/9q
E6ntOaAE/pSdDnwKAbNJrgz7lHw98uQ9/sXrfGU/2EOYfJ+GN5C4PvV3suNyg66hdT+y+1lrG4Ng
GMNrFaoU7kec6NUtTHZ50WElIl00OQPi9u/4Rhl/qyptw8qGETVNef/Vrgqz26LRRDnEzadtIcYO
ahwmm2Nlwtm99J0mhLH8DX+neLmEVPXTokQ4BTkEcE7XhiVH1uuWP7u46tKqwUQje4/jc0JaCCXu
E1PLtItWxHtyT9BeEro7iNH+I9KvnOZ6FEUp2xlYzWRUUxF0IKRqTHYjdwkpEgYdxTXr1IUbVkV2
Rv+5S7X9zwFMgrmIvrfK/KvXQ4T0J3zu6Gwc6qtDMGYuX7rjyBkpcTdI8PAU41LKV/dvrGN+UP/C
58Ck7NwLOpp8aq1ycW0loJnwMuS2xAiDR1yfXp68HomPVAvVAXE786a9bbVh3r0sS3HZgUOyqhmg
90SD17d7bt6m/n+HBf12Z9WWh1sBU67KlntSxa7cLjCTFG/958rWKamLwSRsPFj3fDJwvjMiBYur
f84BGsiRuzRTaQQuwCSYE26e15u3SSiS2PPQU10HVPGxVHXZG9ylMuJucow0lzXJEAteI5TZJHg3
gbw/I9Eh60XOorT5cgAA2nfBqd0mDT98jD2syWwJiZ8n3/rXwMhPMdcT3VOwpZW0RMU5yG1Hgy+3
EDoq0eE2mzxyfUyktxnykvnrOz28B6MF/KXzn6UGDrVlbY48ZpXE6sDPHxlzUj/XReFiVi1Lk3ef
nTsxKpdKefDHVS7RyMD12vqiPkcCFn2VUEdQbXzPBylSxBCLa9nYftyAyVl9CxMKXHPbHG200yof
fapOxJ3cDKFCHRiH8RiqSeZe3T6k/CwqDBANAWmFO8zOXSyJkbgTUbnvTmX6ERvOVdo0OVZFMcYo
BdzTYgYNMPmI2ZVx3Lw5nEUL7IZUXqsg+TO2w1lat1NakoCXJz/Tu7rGROAF5g7xacSWDg+ngdUU
lzVdpWoCCON0f7eLaPjRsn8nUa28rKiS6Y8xIw0sLkZTu9pzYVWiOw9mnbNO1hxyRr9TPekbdv61
UVcRZNKlm2QiNvL1DpUr3DfnzXLSNqyiBLz4/q8vKyg0vouOCiz7T3RpYnaOf2kG838/IAnRoCx/
MGY7HoiUgDGlmshTxWL3Tme8hZbjEqIGZRjsBnuxlELRbUSOowcpH0dcaglTn0iJjks/WIJpIe+b
rjKmVLJl4UGpygcDBUa4UfHWjT1yUOTDvvFFzJihDzmyqtjV/48y4isWVmpLUXXoZFyku3VRBM0d
VwPTFMO+BkktVkm++qe5DngvR1HydPQvp13ofDOn4+l8Ese0SghqNiH1brWXnmR/1JgAJigcbLqH
lqN8eG5DvmS4d5h2anAdFZb6ENUtuh+oK6dzskW0/kdND5Z5rSPXg8iQ46513ez9VG+E2UijCLJU
5Wm7G3yB6jZf9FOFypuX4mxwNsSN3M0wvzgeeCRDC4t1kuy4PSSwc4DbVHfm7qMGzhd50Uq68TyP
OatePVJzWDpiDlRxT85TzW4qu8bmTKte0jJzO+qEldQc6fxAOkQuLGl7lOgcLsy330Sp2gjt5UBC
OlZr+UkUp8fEcZOP6ixZDc/kofuwNa3LATJRYWUbzn5+f4E17rafQFDxJPnsqmLr9Kh23ZnPQHFV
ddVh09FUcjBsX8E4EbqyHcjtJCiY3xFJSZiMNyntaBe3uRhvNnrD7TPSI5g9+QStj2P8A689NYk/
9ZVY/06HXy54c4u1Zq1GYN/8DPSedkjscx8AdgYAoGotQXiLGeej7+9jT2hV+MO6OMW+WO0sDu4B
tV3du0RfACilVaXYFK1oZiU9JK5XNzuOhhPq/3lol+Rys0AwSTDyNDdSiPkJD2YaE6WOrpVXQIv8
Uf8vc+96zY/9xci9n0HaKiGdDJNPTkboue1rBuG9CBLHddu9ualsjzk6F751Xb68+ELOjTMBl93H
x5gxAghtQfYOj5OTsuavpyxSvF0ymUMIzOsxn8T5LHMBHzVBP1XDtHDFNBW5qpYBodjSYYuI89H4
kaCFG4zy88kdQnrIcVvET5bGFYJsvFjOdT5XuKBEFL0OhJKvjnavO6F/94nCTLc8vN/SAmzxp2nX
sWlfqmY9LM4JxbOze/AlvRFIqTqzcE5lN6C8CQpoRZdRKbE5vd+4QwfHWM0X1jF/prnGpGnTNQCC
8RgGENw32LerTRoFxD2v6cFIrAKBjtk0gzIMIWxpkp0OL3Lm9IszgvMxWR9Vw1Q2arAK9XsNeFJW
5d5g8LwvJBpUeEkXJMspJ+dmFV44nme9VcwKgno528TKHZOm3H8VdmtCCA5jhuLg1op27X6HPZZc
CE4KHDa5l0Y2eEb5grqL13/i9d48KQP5NjU24FNrU4JSlcUg9G6yROFwbiLjkoLtkYzc4bsN7jwp
lM2oKR3vAA1gUcKU+FcF9aUOesihnGHoQCwERO8A4KNaZ8RYChRMUo2XoZFG4FHHhY9+isDPVXZI
fS0I93gJA8uzHepnRDfS7oj8xfkFxCjz34lGAfhwuRxfk7u1kK1C1DXS0EFCTqOm/LtVUhkrWtB8
RbsEN7DTSuEHWIc6V7lp36LFQjw6hnf8+XQLGHT5q+YhmwSDDQBTPpIeXMdV0BELwLaOJp3O08KD
CLPINjH8DXSSlyQfYSOuCLssF+ji8Uvzxyi6hkxjAnKquM8jQGLYa/0lRZZhpk4yZrFPwrEd0uNK
zsInF75NaVptbR1SX5RpSMWs18YS2L2j63GtvXh2Eg3a1RRmu7DOp3ETVdKF/I4t6kw3JnUHI12g
fmom1cJFOfiHEPqpa+cCGst9fOZJTp1v9YCCTemH0qr9bRor7LfzjvdhSWOu0qwp9MNaSDodcg1K
a3BbPlHFa1bvZDD8FXx1LJcMbxZJv4sAkR/3dM4cZ6OWIbViONmSuCX2mHL2fTs3Xdr00URFfZpT
h5c7hD8kGRltHgWU6hjxwc2AJ2LXMIZuB1HwAAMlP6ytIDph9KlKwPoeOEAY04rGRGA5DwLTZTZX
kzKuhQ3tdBA7wUUSYmrbCRabSJKBsVyRcyiq17d/xoEuTERbrjPNb18krzK3raaaOZYTr/efhycO
lJCYm45CFl7w5WeMbQjol+NWN6T0kw6A65B6ds3C6So0MJodDOiH6aCba1FVraJMIh/qjJZqFtEz
b5QKwX6AQgR2HsFqXC47e/bFiUak5Segz8q6JCOMmY8fHhQEke5bNMyH2r84KNVNUK1U9DsrFhCo
a38Tw4Vt9o+71KtzqHhLn+pZtn2wTvdpGKxZB1w+Ntql3Zc2TB9sEOdnIpkeS6qOMGBEvVs/fAKR
MV6sNV/0XMDW3UWAW8kGiQ+5my1SWKhf9/bbzv1CCZzX1AjesLZ1CNUdWBgmiIPhrsKxLUnVt0YB
sEYZEK+ySu47wa7vnlWD7Vhn5UtZDNUJ4zsN6w+NnXHah7hmB4Y5PGhsT2WzDa9IZya9bBYpSs+T
0MjVq1QroEWwNkfoiNIc92E4YuZ3KqW1jnWWsaMMnBLqJKcVzYHHjIPv2a+sX4IGkCMMpjmLS9xP
e1P6r5/wVrRWsYwyx1YUWftH7LhCmJj6ySYUl+W78UWc7rSox43nfNbkEoPc+G/IYmkbjqGfkaS4
s1uLdRomwK153m2yuny3SyzgAMgWHpUwFBnfUildnRg7JtLc7TPFhVQmVViaAqOxxnMZzDydsk8g
W5V9pvssN1yEjf8AWo4PKW0bQ+68uiKJdlJOJ2xYsGq5CrqNaHfAh7jLZiBtJz5RGeqNXwZr8qnr
AbGDbVaii/+21wTMaFrGNe9jNqb75URdUOKKZdTiZtiAhi7IloZ4qPYmDKcrZgDeimNJMLlZIbCO
AmUgwboe8EM3K92sBiIq29sghI9npAfXRxEA0HOdb7+Ln6VLVe9Xf/8zRzQ7pj33y8J6BO4n1cL0
HjmB3LQ9Z/WN2P7BXiIuow99xsDAt+ThPC8aB5WZCiY2tSOxF0fuR/vZQCHZI4joDQjDcZoTNfIz
YqOjz+2AAJbxT7lAn9AxlBXMD5B+rScmH9bczm7VJ2XqyrDp4sZkywzE19iSqmsF/Y/96yiRC9Lq
3woNmXaoZ+amdTquAzOOdZ2m5Z6UKkdo1e4Wcmbj+hQlhrRZ1gVKCoGfVvug4D+Qumkjws6eW2nP
aJy665eUJ5AM88n5oXMoshNpsomIgrznJnZ9cEA4ur9l+C8Dr3I297alRoFY5V/OdFhABwv0eHN+
3FHMU7PC4PvV3dIxVdRx1xf3QpLu/9OCwNVmkAwlz2WWKgR+Z1ncncXg/PGLKsckWZQQya6Kxpv7
4Yvp1b1WJVh62rU3xDyi6YclKhpWoK5dDggPbgZeB+wcCEYEULBlRqikuJOti0MwkWWhFNk7LLNS
XPAFcr09TgDg6xV5IsYdc4IbO1kQAETmdqRi+XZx67sHgh6n7l15P691Hgc0DuI4Q1kVhfTabMfJ
98hvZjZXZMZR2dB4iW6uta5CKQVbMENW93k1lxddKfTxDo/qYBQwDTeK9M9QQjm2rHoapSE9CIU9
+DoL74G4WodzOmn+hQYqFWo7Hd+QK9zACVzQiG28RTfqBunMgWoN6L6dtmAmWDWkqbDdPQiTc2X9
VNaiMYbBjWMcMvWJoJDoyECZGTwY4ZcTLjt/oU21hqMTs7VzNgzSBHn65UHL3N7OrcWfFLatjmrG
mZfWLuBUlOj59YpKotKwH4uk8VFboxw8XxrffDcD3sIyjVGf6QG0MR5gxp5ulfOtCn9a4l8OaX5g
P9ZEampdkOH+uyTUOym0mNY7RrCohMGbq7QLaipCPV4uJejJO4TsLnX3sjwjLmOsuC47XR1ZiWzF
z3mNpe4tiLnPKLmIClMMh4mJ36SS0NzwWFFoQzLAF5cajSX0ApP7efaaVEtMy83B2jWUsRrNTUQg
R/eFRZzWeqNU+Fy/YY2hskGAzToCaEWGmsiOWmcqB1WnTn6Jd9EHkgYPbzWu7x9chI+2J8x8eEO+
stI6dCT6dRePzwyAJwo1EAUoSKS4Pg57owDEbx2+XNUA4ZA314dTtl9Eqxryq7DOhfGHWrHPU4L7
9DihzQMuSuwypcjAXWiF53tFYjvh5UcMqleMlt4G5A20hjmGr0RF4rRPgJIhieAVjDKrM2gaKMHQ
zoIISqS/0ySKiBbVpRkW+dEW4449gcDRU/trFLB3g2PkeSsRzu9scxZBS8Rl+JCK5IwwtPwvMmcQ
VGKCb4HVNFvSOGMwqBBLM8bwdnPaIu7rvHUTJA+JGGuQjvUJELPNyew3toI4lf1VHo1FemNsS/Gy
specqVzEcEDwMiS38yhrXL544XylfCWaL8ETNG6+tRM+tbmgMx4GNm8rDu7SRJABjGMWuAb4XP8l
1Ox9PfiK9wnh9E3+CT/jTlX/xEQxDGKH1W+Fb68NpZUTnb4gxxPvIqhZZhFMKvCB0iwPZhSlZZpC
XPmguXmZksedkMMvmyZFxopzIjM7ssOZSg450nBun7BUbrgQ5zUrD9JpjCIfvvuH8T5VS+MbvwMD
frfVtmjXVzFjmutL08jV7ZJx2qat5hR7K7re0NGvryrSdb4dcsWUIFPYL8fSv6h1S6mORGASXhVx
Riws9H/PSPb1V36hfguxdRweH5LRSy2UqLodvJl6CaXAVF6wHGJUwigdlqVigjdVkSo0iZauJV4m
5p0te5nyARJNam34e2WSh6vb/KbpFrVljWVMXeKj7cDYLk+5E0iZIwB5K33OGoSBqOctqv7G0Dw7
WpJkMJozTk9vVKV+y7EPHrtnKsZcLTVvfdgpJEm/CBMgz5ruD+XvbG00X2xXzNbRgtn8n05W2icC
TGwhNagNPo3JAfh5qYkmO7g0KpNK2RF1SohJQm1et+SbOK4NeVV8rsQzU7wjMip9V/SeDujnv3QK
R4Fzi0i9IlGbJ6NCUd44YTTwOFgqrkpAn++bTFWgO4er9Ttr9Y9bHHsKRdHKC4VTZYxpczmvVhOI
GutIdRiz1NywrxpaqjX8c0xqINeRoidhIkvllZZelxAYSnj0yl6MSzP7ZEg+Ek2hhnhtmgsbq9mU
aUl/PoMOs9bWn/LBG1skEJ8rMJb8TbicCOkTK/c++bVGzhpH2QXVMrMOTPRSVWNn+V+Z31GkfJsb
/ErYaNwyxDm5TymLGC/Rjv9utOk544EXIPlHZG3QoZBKze4Yc3sOkIgfvgajopsEUsipMV6WplXc
CzU1N3j07LE7pE5Vclb0e3xZUQ2aGhT8NhR+pskwsMs0VqWkSo0NU68+cWO43AKVHWdoReJpXkXp
03OvOK+ADZ6JxjYb47Zd5eIWukKKF9VC7dEKHES6prcvRFm5cfPbYa935M6DwT/uY2DlRMXWE3Jr
nUfgbf4Xxr/ceQAq8L4BAMWKej5+Ro5zWtb4n0Q/DUdK07jdDRS8b1UQhCk/0JXtMzVo6WxZH9kB
YubLEmGacS7bU6sRiH8WCJDfhvQeJzUR3Z4UR+AXoN6t15mfQcmmdm9AfzEn3wKNQu36qeKRVdLm
6H8wMZXQ9FfaQgMMw5ijvNsO6vjze9hfSAZicFCUvV8v8Q+8xpxXuLXWiiYg4qG8Xrf53x78yAHw
ZbLmIzCcxaBHKnnWfhdILSfC93GKHoxQdBI5UVnSlBjOhH1n4FNtA61uqIjONme/EC8i7myWxDjX
isHAlnEOVX99FpjVdQakU3zIQaEZagV7nlMemA6L4VyukvWPjhp7zh+Ixi7Abw5CMjNkbvslmqC6
Ls+LM17hqSWFhT7L50wbuUl8bfXG33eLvGLnA68CUh3RzypWt5UTD53QxDOKmftDzcExdHhhOK5T
I745bvkr7DU670ffsp0cQx25ZaoK3e7OTSNldU6BCCWvdlCSAvoas8k1WkdLVqnk0eaNYQF3Z9k6
QZsBPOCIitnN9vRM66sLZJvPXFkdpWax07q4Q2SzAzRH87BA4M0s/F8Ro1vLCV0NrTm8Hvs7ApuC
KBkehmJANDQQAr1FsVZ7Vq6h3aU7/svljoc20s1x4KiOUrNiwbWJsfCAjSTOlZ9Gx7bLsDL2VoML
mpeOJL+xfYM6zFUjrsIgElRXlYovekiw9RRHJ/QYK2B0br+zEG6E9L+jn4cBJRhGAPscObPgPAKO
bn0ZLuVqbdEqE6mpfywhWP9CK64Yx8iUb4CiqwX3MpqtTOEcWxUR3+I5IkKJvFAtkA+yVPSzrVfW
8qhCpQ3dgeT3q/RKxUGoBpVPz1kuc61u8OfhWhHC0LZwI8M9gDweJbAvryGJvxeX9fuyD3LcNSBA
HKwsb5CeDHfMt0j7Kz0ABWj1Ek0+615P+9bXpZDinF68JRkEJwzNqiB63M/A0Qoa4QWXkFTBN+qT
AoJVesxDj6D8wCiIU1n04MmWXb5f0csi7OMgNqNy1YfpL2oJS6pDuZ7M69CZfAFHOqI5qD5FAZcu
2ae38Fud8An5qVbtMW+UoiMfXbdOSbQDrUVxRrC6eSzJNp+BokY2nsghRQCzRnplPr4bXeGdgtsh
5o+5iwFIwU+4CdbBPeH5xbdRZEeUSDWYgl6GnVf3+4aTt0pkjajTY8RJpeOhceuhQ6TJQU2ke9NV
aohoaQ1RqJkWyJgXBIMmCcObAnmhLz/YN6jb4A2mlr0QYPm7CV/HB5HTNMzuUUmt64i1w8RgANRE
U1nYWUUbIqC1BVXGF/V7CZZz+GNSIkKsOfHtekgYHawRrb6LY12eh2ipvXUgNLsW6BPqtSGPS7+Z
TcX+9dTexkX4AcNEtZhBJTSdyF4yH/uqrV+FukH/trjOg6XSKCW/SwnbhRa9oCYgLrQKQFuA+FL/
jrWQq0HQ7Azi3KVaZjpeShUKojA6y4cPsyHx/LZuVxN8vVRlDxHvYY/Yj4yUWfMAtj9y1ob4T/c6
0t3O5xyQ3uskBnz2MHUMqWQwJpvszPvHG5f2pwblEBYmQdsqJPTQ8ltY6uImS7aYNPyaTknPUqme
WsglZAnLYRUO5X9+XyFIniT1HeVxmqGt0hcmC7A+BzsfSzBCXAWwWtDLhAIGz/8hBxsm0ntPid4A
+BUPcfj7TjFV47ZFpUeuDY0xA2nArkkcJX+skT6AxnWMqv2Zf967ryWPpeYNAzF73FTwWYzHPMEz
ySbeQAtIvp8nMsrPduOaUTOdOEL4CgxYNLzBGKmD3EfeWNN2Ll7UzDUu86n9Ugy+vFl8Ncg+7ptR
joe1AasuIht5J/lhYcAKkLoWujaa4a8MTqkZ3F9lKC8Grsv6NQgxACTw4Owacsg1Cf0SXYli8xpp
d0xEuipBKNkaAxYqIpJvwyxtDWspKc1mKyXv0vKYwMUt7r6AmY09A/tJVUEpfUoI3g3kmOPV0FP/
CZ3nvmULHfriVYEbeELaOEDgESvNnv21FIz3dh66KsUjBJMNpKSHpgGd9i4SEHaPrICBOW9HxGDo
nnoH/dhTzyR8DhJlng2UA7LiqNBbIEgPjWg1XbW3wEfpf4fMfEzITe7hJSqItJhtgIId+jvEWCkv
WCHxcumcB8S/YJNqH/ek4K8LeayeTkAIxzrl39GDqyXY/0fnkU5kv3Cq3RSgUQ6fZ7USWNV98cdI
a82FWtQUTeOcyZmyr7JwjsBTl1KHh0Lj6USVR6C2QIATYBRZUB3IXc9bzu+29XO5huZbQnuYBUma
J+etdavbgMZ8/dPYbMEtq2sD6kNeR+/LfK/tB0qSimWKThgiDd0D9aT6sbnGqTovs6HUk0ow/XmQ
e8yzYiE0e/hEB5mFgv2s5vI0rkE49EgsdVbbPqeNPaACVVVC1nF/vF9ZfF1nedY803FhHjpuRmOl
nddCnB6hCGAU1eEvoGunkp/gG37UqPkljhuwMnHNGB8dQIKICypOuGP3MjC6ZzgRv9XCByWmKPxI
M7KvEvgqLWd4aQS/w7Mv3azOyfzOAYLjslhrI+KIRkEsWTnVYIlIhJeBawvMGDLBsyPEfR0Xjl3D
VI8nth08+l+6ZzSxAE33T1d025s92oWFzpH2TgQLJyKnwPw8lGLb2zfd8IHT0fiPRuUGoLwmUH7x
5miHHzDV6UCKtT3ngWRSsU4kGfikzhr5lgE0nKhkiZUBbOR88U2OkifH5zbQxb18PW9jzrDTWah/
B7f9Ba9J5ERZnQTAMuf0VACRAdcDik41F/WGofYyWoz2BSRzJBRFuS0cYvJmiJJEmWFBrv24i+cZ
wqNTm7kCZulPc7t4fwCxXiTvp2t0B3NMEfQSKo1vLwtmR8AYxj8lZ4l+1sMhZXnUfwARE4pljILg
mK9grfPpIia+qeUEENxxCXweDs8v/XNtvxn1b1+PRA7gj4584b1TvS7jnIbS6qLPKNJbjZFtOSY2
G0jyiNO4ViH7x6j1m0iH27zeTB+SMz3y1Z6X0c6XtDQYISJ8hL//JvoHh1IaWKJp3TK5FgY0DcN8
GSXsH7g3smlUSTHJh7scp7vodi6/hVSn7twXHHpASNqIt90/WlMrGLq9B+kHUP7IQwAMWijSGsHh
sBxZMEWwgjccuNYjhtAQ1PtH2uclukPnu8ItT3gRWHTDxp5VvTuSGypBJfFpLT4AYHIiXY+DwDFI
nQFebPn1pxx1BMbzen5W99l9nh0771xZv4Gl5Z55xPCAviw34+szKbTTWm2+s+4JoXfffxqx2Cgg
5hi6cSlqWrI2HegLAb6utHee32scESR0norrm8YjmwAUejt8CkU50UAVTmCRxapNAu5hR8W4BXfw
vZS+xMmTcRfrv1aveiitc0xfGV2ONrjOdps+kIfP7liuhsj2H5q8dSBqzJSFt9ULkI7cuSwExbJ4
23g3DJzVoQqEguI31y+CoGHjDatR67V/t5cg8gwXhwj52H9SOo1TwTvLQ5EJdmRn0nz8+vg12XwB
oY6gylYQOfWT6hP2oEqZFNNx4n7FbdTOgOgAdakmGPa4m5tshcQ2XLZVCVOwZthHn122AXy3Vc3d
TqqEnO3D5bPXFxXaf+sJ2kLzFfiU/ZxrSAtWiNsB3HETviGTg3IlphUM/e7uZeF1ykgKkod7eSJt
X8xG/XiU/E0EwgCFsJb0Exg4qrAR+2WLoGQ3LQ3W49HsFQxgtIvgUT0CxDD4QJ7RF/T9JKDtQzAU
FYGlus3HQOVUK/UcxrFN7PDCB/7UfHjke2zauuUT17l6yyuGXesPiW72Jdcu0ESGJdUrr/IBxCaX
FKWLNTaHKwobw+xnTDaDDZv1GrXZP8CrW33HRZ6xmQZkI3QbsvHa9W1tW73AfGOZ98VqE31DS/tR
vUOycNpchGcA8yOW+XGtiPFtxy3PO+2567u+/ICo+jQQR4dIrxLxbWITlJPegYhq9CD2BDgMFp2S
/KK2/lx6+OH41H0727jfGMHXLPt3qGrJqMd6cBkqWotIEsLAHGNegCw5bwMvhM2VV6kVzBEK0slA
shCfvSyvUWgREMizVurVDyTV83GjXyqOIuPy4w1hpNohT78tvLMusHM9hPKPvMgDjFXVHHSo3JRe
eavNqq77J99ssxKtbbyGaoVJFbQjB0/BNqOzwJHy8SobyGNaS254aU1LEn2kzQ7qkEQVtrpi5V3s
2YA+90t3GmtOZx8pZAxFoz6H9HvaEGs7f9p3dQcb2cZnU5DrVJqMrKaFfHGYfSLzUU4ejSWWebPX
h8b7hWz6fTQqWN+qNP3u31jtRPa56+77OiOKXsW/EiKti5udok7IHQZW0FtYIUNjTwKPo25fFrVs
mBcSr1CCFj1kkU9lnp/A+6yqnAOx8sha6FPnHdSnEZM5WbQUu0PaiF1fuTLBK8bHLhqviIO1rZch
SY5IJ931gsG5VA/1ll6O0QsR0t9JVutdZw+62sG3sC9wbQMVUm9QDuOCyys8plqzaC8WzGbeGmO4
5iFjzKi2kHoO4HDl2tYc0xw+EC55/inQirwe9xVPjtgqno5hnyfatHFP0vjt8XbcU/rZKzn6sdS9
fQNVzeu/chfHpEB7ZsKDxYo3WsxwnX9wfiFN1DuGsG3xvBmLZ2Vgtr23Zl95X6dmDxcFVRa9beUy
CjSUmnmw2SEws8CuYgBH4livtiKKJaLC+oTcHG0f7jzphpRFSoD4sgPHt5wCtW/y0oC17meUzGTq
snfYG3KmEo2VlubcN4dXcfWdOvTVz2fo8pk8Axs7ISddCUcJczaG1y1Vl8QQEGCLigqPTVCnbDEG
I/OZmyUJgUQkdioejWNHAs2yFZi6P++7A8KxC/7q2qpd0qWhKbNRmOy7ZlZuQ8ZnUBSC0Wb1OLFN
Jra5biC7PETiAshdp2Y7TiYZJ8gWEl7CCrmn7V9pLtK8GqxdBYlO+a1xG/zB6hgtbeU4VxaBar/m
q9mYGhTmu3RBZGf+JPkvpdaeW8UOit8+2YdzoG7WRKLxhJXdPMBImcrufU2h7+6oQ9yHeyzuhGDW
Vb4zWc4ZjRuP6FaRWHaWBNTWC1W6DQfx5HXVO2VpNoT2CRYgnuIA7DaBsglGg9lVYt4q1xU7UrJi
3DacJ6RAot+tu6uPQdks/TKWRSzIPvZ/LiqXP30JuzOpRDVH1qrUf6IhjPfZv77ONdQSK+0DFZ/e
HTtvdFAqkqQHAYqbaMjV/bace5IgeZkkxY9EHUSvPbM3SgVBWYlTwukK5Az/nvnvN99p9fL72gUj
OuRTYDoic+rXs0cX+LpF/MCnhnZSslf5pLjx+Nlttd/9ken2tvj0sKNcp/zK4F6TD2zrA0Q/sTSi
53hrJwuP+GigpyX2QLblotdKR3WsXK5vOhr8DgsEUMPKdfkJfyK+34tVmXNHlamUYWDWYk1Te1Qk
PEUaS7VSj5btxNKZH2uEu69iTGYXvXjRhuF2NpcDVVawd7J1Ywcik1FIYTc+BlouAdAhoperP3Dn
89iVJtTGeQVO1WuykdJTsPS25MNv+4GA1SAOGtWcuyO4mNlpbVe4lFkbSy2eEwuojLPIMhu58Meh
RcLAwogQ63J2XWQ+bayIzFMS2hAfzEL12fE2yrB/1xWZfXhf/kv7GHctDDN1VNc9UAnpT0SC/bDK
Xd/+P9yg3CyOsRuyZPcqX4d7Uh2ttxsJpgFKmAVSduesWvbOS8LlrbD6ZNz6osBE7qfQ47Av2hhF
2bADv0qQWIXH7beLUGY3NUeuqcYrXRyNaO4icq9T0/G3MaMoNMjWGHbeT0Ithb4l4ljJEoNSdy7K
0VN5VpBteYBYnfEey2jo6mTUjDb9RmqYGvzgDwutpFRmiTpWnpkWDGyW1Tzl6wnCRqrK/QUdcIVG
ONPuN88f+RF0Jk8L/12ZnyQfjETRRzMKCfU0lbEbYVO44+XGyEUgE2/tZAtcYamQyEbZjxIYYmpH
Gwgd3gq/8C5v2nRtUCdWqhgpsZ//jq6o90muVqPDUljq9cgLyBSYs3nEYS6Ue96QDF2OEAmN/9w2
C027vr1lMrYNIt5k2uswnz+rqXGWadi5VN/a7SNjsx7Y41Yg1IrA+QF3FVegLEauEq8uwKF4DwD0
/NRVAnnX5awfbk32o1Lnn6wZTbbqgIVkKkgYL+nVtYkODB7pegXLB1ZQflxhQXdcpC+HnrTi5N1D
HmqWWzZnrw7sm6pGaA6mT21gB2iLMoHYAW0wfSPhMmrCctELwiPBnl0OeZia72MXyHY5pyjHaGkD
Rf6y4I71WGYMOX2X4ZTs9nBhZjPDTc4PErml7p+wm2S/T3s3m4AXisUgD24S+wAVkVzT9KVr2/Hj
LAtSmCbR5JyBY1WMwoy6Loqq3ZY6I4YnoUeVzTtUpmv3oTcDOkhf7syPCdMEUjmQ9vbKlTeXecYX
7dlVaLJ7GimJ7gHLpjUuPtBXWwxgUl1EmMX1eJBiDeANwcZ69lJAKSM0uda6Oe9/3RPx95WSJZS9
GtSlVVePTPWh0J2hRYxeDJhT2HnKmdIUNMTpPW1ttAj8KHGh/cxy0K1EyV5IFMBFRxCSIO2Q8cxb
bwjYSw0IbEf72AQtbdmpDSQQUEN9CZoyGEL1KoeCO+5bVqwrZLgW6g8ogf+Lz8jR/Y00t6cjPjl9
N0dgR6nGQeRvvrSaFfnt70OafH1zzAhpApysG3ioJbzNA2Yqnk+IfwY4pPkiAqLJ6Ruup4ljukWZ
etDpgiNY4wl4YIPPqj7SFbUxti5lTtTMyWyFAJhRZBUnqyPjeaO4og27k+btwl00YtaEmZHNW7Za
MoEsQINGm5xjX9wz/2QGRCloFSH8EZHx3Miasdy5UsAimHrlMF/N5a8npp7JslHV9SHEg5sgKRkV
eStW3Tq2Dzze775YpkGcSvDPzwvBnpqbPZxYS0RJJifFkKUqIFeaUGOVpUyGOvPsCbEKtI6iyf5P
Qz2ZE6b0uCxgyFSbesXpvCBK8Qekto7J34D8R2ddAPM+aLnPCZPgbeDxwN1bmXy0Yce8tU8RvMpE
2lVhwY3P5UxWKLfJ9dbdi6Aq51rM1bY+VohxV+rlsgieQJrAICmn9BnswzKmVGRcbMi8zoXVQ3hn
z9yNAajTr97BL8AWJBr97kVWV0lPyK1qeYj5NyePZIoXU1QXkWjB6uZsxgZZHjinYIQDTgfDbnQj
wsgSIxF7cC6h3HUXS9ni9gTtC9vSp9Q6an8k66w7M44YqgMv+ORxlpmxsoHtJgCtkzJ05bB3GnT0
89eZEERrEeTJxGIbhv6WPHWNbyOupbXrikiI0IC/JKbQzo401DX3n2r/xHp5khuQQv8cUGrQx4mn
T6ABsK4pkezVsfk6AD8Zk7qs+2RO4NNuAyCZ0kkaVjYyRkz+rUHbywLqz6FGnRYdmP+WxXmDk9aq
lgNGWtF9Q/VpiRU9RsOUTOtmqadyaY6XUMKODbtZ3KF13C5XIqAQjQq+QXJ4enh3x4Dj3IpkOmRJ
lh3Z4QvHZmAVmN78lni+Q2t/fNBRE1VzQc5SEtaUdtWASFrZqv/lF1OfgtcnlnYuuhurlRlhGv+s
q1S4zW0qEjV0+AwNi+OVQ45cj6kHp6lZtE5uWBL+yOqE+m6n6p9jhBmUs3NZ3Bc822pVav3CUhwI
+IRvMURe2dCL41Q3GF/M1NpRFs40qMUJcMGwmMCEquM4jb2Rt1l38vLAjp16TSEEJsW2BpeEULMf
t9qNwjqY65sq1qTpSTWwmjSh2Gpr+KtnKaCC7wos3EfUozbpCfRbnMXbpJc3adVPumo90WF1UNL/
LdIw3JaF5mTnqhqBCkw+rfMuUVNNY8IBSt0YqPMVS1K1e5jHUKWpi8cejS7tuiQe9tu0rRErLLaM
4uPeLMO14W3JBANFtdlgfiH12sCQYsHgh7t2xmTXqzbkHeyWXqyuZ8W554acfyAQbLyn8oME3eOe
RFiLey9cZfBdMJu8SxPNx89ZBcihXAK6ZEgLsXvE6Z3va92P1hLNZUhSr9XE4+8AGIBVrWrv8j8q
yhRVQ0iUqmSSKQ3T7iNvAVEYFRL5s1IQQe9c+diCpXZ6EKgJBsRvyXJMyvlQuMnDPIKZMFzT/8OU
zJXepjyciDXUwnD46ODj6gfhzV8m4azCcmoVKlCwO6mLdiel423MDCDdt/o7xVIF4kppQpkLMklW
cYj9zML58jGmqlEVbNuuD8IyiXz6Cj97kN6m2WjFCbkE/cUIAdFkmyNJyRXDrtb7aHyg3kx693oe
JrNO+8mBw+deW8Dc9GhNLW2d965tvVA0PJgOMXB2yfXuFrDfkpwfU2LPoSTjdZihbkuCG7Ed5fsy
hPAAGSXh6RI6nTEej86QCDxQbPFhNWpuDXzWkqQjesOLMfi848DpU+pEOWblTtvZ/r8aWSSytf1b
lRg2Pwd8i1GJ3R7q53dD6Jwg2bPb2UwBOkqRhlzPk2XY+R6uBLc4TJclI5TBkAKJXfmlmABwHtFg
XiscxaWI6KXks7SdoMfN600kr2154xZMLfEwAWniTR6Xly9ZRuQoAtWsEO6/3ounhVdxgd7zfE0x
M8B+6RxMn0g5ls4vzBmeWqgzXUS4LyRCI+Sf+mH5Vfdfncq3DzO/OnO4EdZWvMOoGMvLvyPRa1n0
At9WXfY5sjg4fUKgqoLzwVBx9UOevNEooGUGuX+bFX/UBwHhEclc3WxDEpBp14SkfaLjQW7Tajxy
gucJwDXOw+V4Y3fIvb/JH6TOeoOqVJ3ti1jtYGmKr4DpSBpPqAsvXJH03pgfp1N4YCrbMrPxlERa
myHplvll9CuvMskPJBb48p0f9zKB1J1VhMPWln4ouFgdacBNvVvui+Qc33JYe0HZTBzaaVRAhAqB
wur9LLoXx4r0v2l1deXgyAaDVqr174AUKSeG8a0gEnnIBkMxyIChYxjZm+wJDGuHrj5RZHRR9Geo
c5wKOnG5cUaorLsPXbqog4b6pcBYCa4OsJ7/QKSWPrtPMLAEdif/7nJxYWeSz9cc05yIVcH/O4bN
hh3ldNNfbTKlOIlS2SAeL5XQdhkaadYr0Og0ju+3vkDYF0bCLazxBovMh0O8D1ocy3BJ7u9iK4LE
RfbYxqhq/eV8wddOOleKtfDJ/ybJSstrlsMC0iZ2XxpztaVfzdg4bBEsidzXQjswCLYoc6N1CbSG
2Z/xL/opikyNzeGm/XGrcp1253JFHfhUiVS6uHOk/w9rbWNlvZPHz1JTzOJoOW2kgNIvhUQHSuV+
BB4zt8Nj4Qvn8tmWy2ib0R6khhZr1csqrrJKmvmW9Xx9cyZ+Kh2NMlvfHHQg4PP3NKxFBr9KMdyW
D8G3vr8M4CSDcSq/cgOQfzy//6sskfvc7Hzqw3ZFvrl7h0lwYhN+Ekui51WbwHjsUWlJk7MipvZe
Use1KIGkxKvpRIrVdGXh5yLcpip8eSmKh1fa4z+lCXK2ta23qIJZpfvFwTMPQQuu/wfBQzOaXrTf
hIDJiwkbuTsojhoHOqtIcQ5vsevUJZRMLn0/14YbDJWldd6tgyA9N4Orks9p3h2mpUslho1iiaOs
q3qgz4B3WIR6BaCAlzHVmXdGnbb3NmBpxYhiRqtsd9PAXuTfkd5aMIb9cWK7WJnigX72jadmGkwe
6Z0uz8MS7wAtLC7Qsp2D/7k/boWCpVjkI5aq5XMn6cXqM3PvW6k67NT0S0f9S7u7kbdTthZXt3WL
3DuiPUjmn6MhWWqsjFnuyKIsSGF/dn7sa6bXVG0BY7oosiabvGsJPArcmrHCJXpR4oLhW51qom1U
1UJN3UUscFxnuL29kxwStXqYgbkwEKofn4TwEL07lxv91WIREaS3rGTD3996stgzgszvSokhJ3r0
yA+7ZbH1IJFk6pKS33MMwrnjtZ9VzwOQD3srYM0Kg5nVRY1RZKVfkn4cAUN07srJgWg8KQDSj2w6
bH6Xzm85aXT0/3q1C31plg1Y3rAdTsQyLZV/pLPzNN1In/0TwNEXYapDO2+DCuPgtMmjeZXv2INS
03jX9m/B82tzhicHmw4EA4GCTjN8+Pc1glcPKz6zliA3Xv7rJbaVXDjWlRWUfWo0w5eEKeXcRH6n
MPZ+9g2oKIDVWKYGC6ci19zdgpcI/YEzuv/zP9uC4PLwmot6ZUO+Zzf3yDsvcJ87uRWRaffY/DQf
G50eOycSRKH4VI/rrfCpfS44cpQJPcWPF195rv/81idxiR16fTMEMSViI20HwtlTUknYd1hA99H/
9YWAHO55UuxBVuOIGcY2xY8Aur6C0xJhPlbqvZzY2Yaab9rFb9u+CoaldtEy/W0zYtF0wJ27ikst
AaGr1r0/iEaLwPi7IflBIEi49q0EmbxNONy3KkoNxgp4tWFfbL+kbaylXppNI0+etAQ6FjzmAV1a
TA/ichzcMeDJj7KWpPRA3N0OS/Vl/iDOVEPBOmyw9L/6LST3FnAsNiEKC/dkD4KPpJFL23Pscezp
r3tM16ad8kkJ9t2M9vQX3QK7J2jALlZF+GQuDEyZqofzH+65zAiPKA3d2cNPiutRr7rAmSir0USX
e+jgiXWKu2b2eRGgoo9jnJ1gwZA+QY09/I4BwrVmzsiMaGlLXmEsfPzDmyjH0ioSubXUIVl+dvCE
QSvDETf0Ti4/kbuP/ShiAzMfPkeloSrQUqzl7PfDZ0tS7Uc/Xn3pEyhSGinfTj03ZYhm+jLp8qaF
eRcU9ddUMdPoyDUUyze5XFd5Q1t5gEoR58ukzxWtHOn2uCuqgj8CEEgzI3NDFzzSBdXSrhOTAeOu
XqPfnk79naCwHvJuaexACH9W0uMxhvy8ZD/wtL8o32sludm28LZ64uA4ycoPi6osoJR4KcLH8bxw
LG3ARD78/DrWBs+h5gxidEosMsBAckuDG5YXzqqIj7sTdKBPff9WNLkQFRlzQsbBQDb1fK53umOM
M18dzk7vKP/pXCMrQyNBM5yH3vD2yZMl/3nDJ7/vjF/w0KqWyI8p1LWs1yYJRGsmnbNzCbtKbGP/
CnNo4XUWJ33gDb18VT4d/gmjpcYPVAuyghnQA7ZMpjh5q4CTZBrOLg1QmYAtLRqxcSADXbOnKYA+
qJGJL6bjtE6a1iiAIKfCXSsNqpLL2Uk89qi1p3vsX5hbuD4auBgdfvw+h2xf/ricd4g5pdg0YtBE
+hmiYAfR6+w6FUKhoiXomNRJbKnc7XPI05OJFxgkn08EHnMGbaOduWFx4GMJxh870A7nykmDSJPN
Wyiwn5WEkIF4rMeA3R9gAUXEZAoJUsIv6ahbL4Y9jVX/cuN8VaD30lobNyucG/sRhoFPm48pxXyA
lHOycM8t31axrVDV2hhkSDF5zqUUAtg8FFJ1gU4WvYbf3rC/NZx+Op2CtQe8TPS/mm2sBk4P3uLr
2ND5Nr3Ifi8IwP/gbzXilGlO4I2lwjcwIDMpkizNpR6puop/vkdzYgRVYWeXE7R/26mzl6Me90Hr
iI6bF0cExQJ7Bj0cnmxQJyAngJkNZ2zTiL5jSUqlGqN4l0BLTmaDtRVK2X2CKvUb9hm3aJrVu+NQ
NzTxExMNwkmCsKZUpqdQXnrjtt3xLCokN1QNs9q6q+vbE+jxZ1raLojgfEzL9HVUyNk4YDXXBXr+
PPxaUs98CRu+clr2qVpWqmR0rvER4R7lVfLFr3oSyX+9Mg1gEU7wzQYSpUHA9ZiE02FuUjRtnqj9
MUvKbamXoB/6iBKAMYYWt5/WAhddrMji8OlvmL5N31sPZTzGzZQx+trFrWqFR31WaZt25ypZI0sY
RVTDSWh1DspcB1H995umaDAFfH+t5swWaYfV+2gC09Y0v+aN0/uJQqRzuUzrAkHUYp0zM2AE++X4
qGMrh0JZTAgu8FRjoG5YVSQph0U8BOoOu3vee0ngRVcoh871qxmnzpP2PufuR9qfxNlxROY52w34
YJ+R9MLjv+kCPlkI2C+54IzqHnEyjd3sIKEWlrz9BLn/PGiCxbRIfi06V1uiwW1s5RRRTq0XYA0y
eHy0wkDqnkqcKmHU6T2djvCc8vVKr1jI3KtDmfokDYzEJg/BDCp9L+1E70pYu+PNqSNkXn6YmgAQ
EHouo1XuQeE/qx4g5BNOxVh4loe49W3wnspK2stRjODCh8Wp/qE62EIRZvg/2sG6wHDkNutjc2Em
rNzJaMDbCkwfr+RPEQ37auKQ41q7bpxzYjB9TQ97c32f0ZMo7Gx4W8OT9Za5s4X5YpgFywR4xYWp
RG07J0nRWUDpgBXQXlb+8jBK5hEuN6/zRxEE6VmqCSlyxe368D+SJiCLN9Oi6ZHfrYE6Bs/174n7
om6sFos8CKqnWsVNIWyGSIsPS83+LtTXn4Bj79ThJPBDksvsxQqrZPT6k4K4C9DbbThJCsy5N99q
RRu+xG7j2CaCpvilN7OJC49rzjrhKcsIIiy5UB3dmikr72/wSrXhJp+yG7/Vs9CxTYqrsS3nvVs9
wbk+1mD80fcrBmqzSThsvnH4JW+1Ertvsk+E/R1OKXgMxAJYU4ywSiW+3xfo94v8f6M3k3IREPlP
jheVqpzgPEMXSyPVMqrXUlzDVvnWgtgyNdIKf8Y+KXUK27fX3slVPWqr/ksM/akyzdLG6/bF9Mp5
nomcmPezF8d8W8R7kuMVTRtABEr+QUjacpjdjC/4p20xu8v9bQEL+HeABy34zTNtn01aMtGH+YY2
nSjXpBmdlT6iEZXhUcRg/OVtsgkDaAeEQ8nD6cEgvFccKKMFm9YtfeYmsDXO+7VZ4R5UK9DuCBTg
9mFCW8HzEFwNk/95LdCIKrzCyOMUxPLkNhgoCM54rck4WI7yvc9U66Txxnqw/2i/4qgxCw+pGXFu
XhEwSFqkJqcKr0IJgILkAstFOUzPwejusqbfaFnH4i700dK+qov94DkHU4mQEV50SVW73YPZxKc2
heGUbMuj8g2ffVVtjduRHxMKmS64Z1ZTPdpaobIVdfsuQBwwqpTRnjS7Vssrbuf49V93B1pj8lZ1
ICLl9XagCNFxvXT9z0CPVt3wiDMrxKtvZHKV8/OWiwPIlWVvq+UShMxA1sQrjoPsda3kxMcXu2tH
y3JZC7zAbSfsIRnKq16ghHyhdhIJ6eFY71kb6nVffIDIhp0JfL2lB863/2w69O7Ed4BZybq+AlfU
m8fBjaI1rWTbHxb5g+Zz6C8+DLIi5dxq2lKr6j8Mkuc/jP0VYj8kEL455D5Tynzj3gP4svSTvRDE
JQvm6khTmCbunnIF9Ih/b0TYjPMLOOZ98mWnFFAVP0XQABgtTsWqmqQqciS5tyLFbwzNd3JDP+p/
AIDNmLPz0vEBXR51ALsZpKiFnnkdq1kZYvqO2LAD2rC5dp+sh922bZvCr31moeBP4GbBeEB3Wldm
TDmioL64CLRrsz4HEGud4NmcbH6zz61YPdVVHN45Ivysh1LjdtcbDBcURVHhqnOEb4dTH4lv5/sm
gz1WZcwvCX6XYMAWSZpECdS1VECzUw97nKONKvj5bYZmb/ebcjYAAe8Pvn4OIc/jSSeTXKIirwUg
UcfP0GSqUVTdVZeaDWMndDHvPfYKLm0zEllTvQYasGh3m+rafePK/c7J+29au0Ut8DdMPhJdLHpT
W3T0S5ORL+ivOygrdEHXS6DDsP7ZAnOpshz0HDVayD/hY8FKPAYWO7p0MO8k7gLoGCm1aAjzbILS
JxQzGlyinhgJgQzLUVBtC/kBNgFgs+xJ4DAT0oh89oevHuBrFE8BICQnvl4CzYzLGbuPi798Jwhq
jY+vJD+qPGRjjMaIlIyY3INIjI8JbKF1yI+6MKa2xSsB+NoxuGLOiOuNV/GUPKq39D6s9lc5GD0o
xWunhlDettvPoE+UyCJ0CH4ou2lC0iXVmirQEaOQZix68WpgFrZ2XmEII/nuoVPudlKvVp1XsimL
1g4ug6Osxs6EdnQiPwzsCn/8KC8AI6nf21cYk4bDHI97ZIxZ4MPVxbA9/gJXfaGxbEn0/kq52rQC
VuQ6xZ69538S56trh22UVh6NcMMWVWssQrl8fE7mVnDFBoJgpFW9gCNIDqEZVDkZSue07jmw8eyG
0x50AK6bLxaFj8rRHQ6ztipTeArkF0IHCBjnZa4hyj/NFPHg/XCeyIhUwDRuIrhRr1QZj8sBXNI0
FMCZC5FtAbXvkKVOluTvZJI58IhBveFBG+IqkP7w2oDNYvkdHa3NNK3JZIcTl1yYAVipFz9qlst/
gKgU4WQjkVnLzpeZcK9dIueXM+ienFyypeeenZav5cV3VP3DMOsAgePKJkwlvXvKzY38K19VKeTn
DP+KgyQjiEzI9ToAPbe3H62LtCU+6xa7l47IcAgenQNzeNkqxHPLM4YuGVg5IS++v39JYsRfHFnc
2/100SKv/i7xHkRTpvXION0fZ8w/D5pTeLz3Ddp7+Vr3erf+yzB8Hqm4+NoenO3hvmPYBdMGF3rv
m4RG/0AYtcqu/x9FXrTct+akGqQkWwW05Z8YfhRPigXmxrfEkdq3mvSfPE7gCgxZy7HPOkccRIq+
PwciUz9Zgo4XEIu0k9vUCSIiJklqpzajYT7EMtM2WRo6AJjViLOK2f84dyMoDNevp2bgzuSyDCy4
Swvw3CffOj4XEelLjNZ2M9gAvQq6wkTSONejs8p3ByJGLOmvf2LuSVgnIOBRAe5FmVBmIJntrdt5
BjmNNyhhci3ABywQTF6wP1ULAUHzLOe4XOZWywlhmQc3hIqqVkfb2nbrQyLcHDigMejWBpcAHPpd
1enUFSrjZIDKk+OxzUlNnzYa/QbaYKMilKqlIgT4FTJd8z8Zgm8W2gc4w9k+Fw1Z5chUjB1vURqc
t4M5qRGfyYHzr18SpCL/QPr/83c2V/f3On9XoEYqOn9YHlQcHmNzkRcqoJvHOIFaXzCqr1YyGqyW
7aOM5+pPLeb3YgAk7Pnzbrp6rKdkp8cpO6Zlp4xgaVHcRBWDPgEnPq73Gmhq0CoY1Nb/1NntPpV0
iV/GHrFw/hwtSrLqO2MbFJQ1VcRdQ2nkWOVEyjwku59qUR2zOp9CsfFen8MJcnVoBI8vrjHMmWuT
x+achjJiFRM+GLVvm3tY7qNB3E0A/QD3w+oL6SzjmyU+ftWJlb/MNehNvczCU9lyhrzLoL4bkHKt
rd2qyOjaXtt3KLKVvK67/SlMrZzVqnAabOr4l4a7Wq1C+SNRol+0iNWUgoKOtxzjkWtvTxsslFlx
ca+suGMAqYXwQ2YOTpUg1fB+NRxF4xdDT5L/MdoG5RbeZ4z78MZbsXKAz5YfZQgSCVtwkB7XubfI
QAchyxejcr8mdQHYjaR3ZQr/+TLf3T8+1bOKlCmcvorBWU/vj8My2zMp7hKfsiAgHWmorXJCQcdS
KEXoPWvUsP+lDQ5ztgkvqohnoF2tHD9BZkGoiBK7xHaa4SA7cmkCUSerkqIBVSZfKz2H0yPG1RUo
x4lxtPyiVRu4V2h0z27jNZKE41ec0aEUcAsE2jiTY162InbVmOamwhQDQiZq3GtfS0dTxrqLC6Q4
Dnr15/ItGQdeTOQyVKO1CwlUs37hreOqrFNJqekQsTW4Qj3/wAfTDcNCSRCkpXO4GWwlbporCqXS
GJaRs1VOjEbfVSgI0XGRHGn6eqjSjEqugutB2xSMIDIl3H6yvRzIZtBytpBzSNpP8stK14AJ/UWv
S2QBhEYHUZZJqi5tu/aOHxSkgvBPftTGhzwxOFPEyyqYvh3g0JXL8/3MAaxoxOAmA9aXLzhsH2Yr
Z3rspKxI2F0Il8UJyySCgzsPL0pCBcuYOfl6G0pMedC9Y6Dv5/bVsF8wi24IZHddOm4UISxIK284
vbyT5YVOJGqHdlOP0slSmQY7nlS/No9BfnuM92NfYWB3cUSNMbPWGSmzTqr9ynEKv69jZ6vseewt
4/7/or8fn7YrZnNk0DM/1weJms4ae+t867sylYe2+i7D1fUaNDRvUEkkOyO2SK1frYXVZEbgvcVC
MThFz/f0paYQACEJPt51vfGQPW+altt1AWuyhXoXQW2ymP2kzZeiARQFDKmLf5I26ye3HoU7HESf
y2hS9KtTnK56vnSmaUC/3p6aa1jrWgWa1qxZD+M41TXyA/aD1Ci6tTWG7KI2G/4NEBxLWu4qQmjK
hVgD3BRviXg6oPOsdX3y/lobwfPOtUl/y0jgf4D0wxgcM2PttHGn943JrsThH429QcpcRqmBMCni
ZyiadfKRXNjqI9hUJDfta4BZc7yDNmP1uLuXJooe+hgeK36U43oGXVbIFoVbc+EBezqskStzhNZZ
phMK0fYOQtqgFOczvvar2PRY0LQ95bJ3976Wr/bU32N15/Hf9Cbsurc8eLawkCWM1CU0LEsnHraX
p/jsJatCT8nMa7uUvctXULFG8ukYqXpGVYEqeBuCDEoVpAtWWTnvE7paqx3ZmLy3OHu8oRFwZxuu
SySMZtvsN2h9jxV3RzSXV9a5F+W1v3m3oUnrEwniP0ezIxw4UUjBWAJXyYcy+7nUrZZe/9PU9lsE
a/3FxfThYGtrErKYzOgFbcc/qb0V+pGilPRFEPoBKrmCHeRa+MzxjCq2o/y76f+rNBOMB5kUFcoG
NfeG6Afx3aSOYTw8ykMeo+O2Y212Ov4NonQBUFfQVgU9qEdt23/Y7KI7LQ2j4pvv7S2Xq3IL4fX9
eOgOkOiRrcn+V4uKt6GIXwVnUEKituHp8X2em7Av7teKH7DU/mIHegIOqiP3gg2ecOdzvTdwEdf6
O9NihKW3czLF43Vm4pXM/E10PcpMtW55OtauLSazA8MHw3bFRCTW5kebttdxDR6w0oekqcVW0VKW
4M012VklnN9ISl5ZJs02RvTDIp3kpKXdAyZ1zW3vE7dKVd+Pif3Ls4tN2zAVl1fJlN745iHUTYzR
cQ6B2k34rKXXCJ1TFte2uCAAxpKgV4lQvnpdK5u2N+b26cb7JMtPDxDD9VPudbCog0NhenDesVS5
wGXhE17mgFlYhUqiAucxfaFV2bodC1Wf12f6pCoHqHtJMWLqI1tAX46sBL5P+Ov6xdln3gteP8Yu
0MVgIUbkjzxpzKPIHMDNzxFXTReAXTq962kBFICliWHbcB04FWFQ44Gt1iDxe3ET6jt5IUyDVMxB
XBUW3GdV9+h5EG9e0YwnGK2JHrEYS40AZI3druiAfOcQ8SXkEfraGZhlnjxdY2jU2POOz2odXu5f
Y43Y/B7YDgc5twP2OZX3BzBKL7uJGb4NgThuGntTOt0jeWIEKtEGKL+ruOTGx2bIRBt8hq3ECFd1
1Z9kvd4wmJ2PhEwm4vZZwphKnIEQxXRjg4HCjyM6YdAuDt2yauGHw/2pzvUuY807oGR5x8f/M8Gb
mK11RIRIpbCHa5f7JrCFF/4TVwkQ2GcXrgTrIdcjmQSJN7UgBBiXu0y2hrd3pceQsszrIc/w7A64
kK8VGrExNMZ1jngBTH09EW2sEeOg7cH2uT4UjhWmfFqxSWw7owGBE2uPvxEwNarDZrG+TxL3BabR
1w4Y7qmaRE1pW2cN4lzK9hvjdS+r1jvuZPPCUUsYSk+7wGrb+MuGW6/Ux07lM7YHUYlcfqZD0qP1
bg3Jw4dQIN5WrxA8gQ2ZpeP/cMYYbJ772KTX+GfrStrMYbJts5CI7yS8BAAtB4rhr247PQH9Q4T7
Odii5O1bthOWazDhikiPmY4IaCE/KPG2IJZ0gaTppe/nefuPl1FRRoUiKSNZa07HRqdQKrJVdk4W
i3GeVK/AuRtrqKvlSkVQSmW+u8Cnax5i1cK/Klo1OhxKFtLZjKipN8T7c65C4gy6rtVuwYi84gRa
WRPKA8e6vEbL50Mk2KVIhViVMLgjd78/H+PYgm9zsMjxB03yC3rkfcoOpb2fFsBsdwCaDvDgqGe0
IDw15/fE1u/gcFF7sfuC4lSH8R9ATxUWcbJ39WkyBZtmgkezoGQbnDv7xeaRU8p3fB5TSJmnAan7
raBAwY03Hy/7rWYx7G7EzZow83t0cKywRPwqv++zJ97/Z3B3iW7lENMVyC6OSOcCLbEPESWCR2ws
JIS9ieQFLcPTRbAG+w0jT1uBt9/5RzdfOBTMVftc2V09I8kQkzeFzqvPCtfIgyorPqRl9TZTQagX
4LBB9ZHyl8ZGNXKnyJ8m+GsC2QnH6pLV+qSlOy/5mm1prY9luY45YeQud4KIT4NB/u24nPRbdDO7
5dGbQGmuvyNcrMa/lpr1qo9/j4syRRty6hTWL3jumNjD1OHzlJGOOQlDaGfkZUiE/bruOZ60PpoA
foh/3UK8Bhlw2PuV4sCnOMR9T0JVyW/0aNSX9BeuCMQExzeKQr6YuDi1WtcJ5lZXMSCBq5mLJBk+
PK3jSmlRIHuvf0AbGs9qnQfWAJz557AfMb+CL/tMYt2msUngSL/crgW6kedIC9FNMQJnIBHIsPis
OUPYn/4XouAIjVwLm0qJnBrUMQIwtHDUIyuXayFuf9D8yEiIiBAQSWg5wtXg9fyzOqlJfX+FbbNQ
DmjHsdctoBzRoD14B0SyGHqczK9gVP8fIK8NbdmzUiFISZ08EE9zonG+H2vjOawHCOHk3HgyeRPg
LzfmVY0fzq+NkAc2stch/GsZjta4StSEnxgKAm+SmozYYhPMLmq6jXmklnUUzMkpzl6N/rdKTGSo
/QzELrZyT8t5IthVG0ZOEVoKqCnQxUuslqEQOv+/xiAHhpaH6rJubDc/n1BmnKV4aOv44uF5atcL
YpbKnvlRcvzVlt1UWXPb5PypxxGZ0kbJ/J49XFXvZlqeUKirhwKeAOuDl1NJFm9xjR7PNi4At4iU
37Y5viAG5ZAORIjzFVDGk6yZsbP9Td/4kLXwSQR+VUIh7ZcSt/tZh+sHUfXQESGKU89DNN/3vZeZ
r1OgSsxrk8q4boGPCK6M83ausNaRzi7WblemObDYqQWYb61i7Yru+gbU5ADH4CMp+W04FR9lxe3J
G62pi3NM277AdFjeOmN8hHrnKADqwFzx5YaRwS1hkGmkec3MUf8A19SmmATbGuLZdUwMIy0/COYO
GDntAAUEIoemAyu5xXK1DZ2SGTjaqcPyRn+EcUApnliGt6y9FYdGQkpjbUvatKgbqkawuss7OFGx
yLBaVFalBi4BFI4d5HA371wqUMfqgaYv065fLza9m41Zi8nt4RLARg5nZaB3TxTnykWv/3T+6ENB
UpJ5LwnKDAZSRd+u+Pl7SXTPHwYRoDXN92OxQbABXu4wtghWxAoXEzmBnZtN19O0Ir8jXv6rfSu1
tIPYLNzCnhcV11FaWmQMO9q1g60Q+kEIFvZtgByAQcGA3jAcrRlhkSqQsHKVWNXq9tZeiZoclAmh
+TvCEe/DgOAWFQLQX+gmgkkYIuS6YlQFYrYi2V205+/i809QHzZFx6TyAtbzCOTj6c+SAYa5PLBY
8HTX2KuzXnvkPwjRxf7wqawOaeXWX530KFQLslgoS0oHsMOWD9mrArR1wAqheMpoSA0QZYjAih0s
VEcBfUOy/IfDJImGN8CBZJ7MynOgt0XbMGctY+Mak6bLn9nEbrxbx+4qIawCvA3pUKsKWBSz9wO9
5NlPOO8xFFjdf+mHuw+9rS+y+0zxcjsB8yxPRgpdgshkXPMHCL8zG51I/qt5xtumTR3gPdpE4QPr
I6TqMKd6Oq3sxqy8wcB1MuOPjKJTNGsvYK4HzNUSK2nNNqSWevUf4hJsWAjkafuaPJOdbeu8RapW
+mTc2b6RNyvBTj2qkpO1pr9mW9w1awLx3VXf04mPzmKGpSVaHx5wL4kZM0rJmNxpfbGs8hmxKCcQ
mUHCb+jl9uoROgpxs02JcgHkPrV3g3eDNa4zIK5o6xjFQOohDtr0GtFfAXWqcn2MIpx+i3LQ72iC
XsviLC4R9Z85GQbOU6CRDJDM8VGWRt9l4HgqI0g5bLAp/TWgNjOHgkg/BzxgJtGw4Gh6+UJxHXr8
7520FVHSIMKUv+xedYJQAnfi8++Qp5RRE5h/2VCieOTtcNkm1US0K/Ebyga0eUeAaIw/iY+LJRcH
rSH6TgwC5F1GP6wmksNrVS3ZHlOyQHSnOTcfF9Vzke/IsQWV1q9UZSdL2ZHD45/6stCSrWnfxUCC
OgrNjN2n4Pfc8pJLULlBge7n0fsHfY/IhNgoahm66RMn6KlqYBdznttSDJDx9/ie0AnGu5J3GFQK
fZVJKb9Q2yUlW91CRMzRzGlW3n7wlxnZN7DsnuUWhNNV77axmmPhzCBbwRpTLVb9i8jZr0e0Km9V
9TjCsWGGBWCHz3ZZm122Gz1kG3+Q3tCxINZkCAktAvW6juLESo8q4e2n5oh/wT2uvE5B2++j2xTt
u1wJQ92GNoRh9lgcUjW9rA+HNso0AHMqoxjWF5ajNGlPqfPbIOlaDaHInpnOS0fCbXHptwrjFIox
ZveSvERnTsqnNJClbcLaExj3V6yUAxjB0V/AfqUlA/jLSAI8m4/wPBqZ0f+YhRl7xPgjdrSIWlB2
QviH7v1evjoUXJKMotsBDR1kwnJexN6fFHF6VvBp0G0CtS7KiYiiGIn4duYwnzUFjKUxuZl/Wo0e
QgvZBOBgMO0N08t86XGa0PMTSjPzwFtvOQluhhzDMJHw10INpYmTBKR+YwdIrOZdRhSrUJyEVja0
oB51s+eaxAXsiCfiAsN+cMrsmj3q6sKq40RJ9sHFCeCQz7VvPbfXTjU7kSOZ83Sj5J7Vu0V9n44v
R/+CPaNP9HDJ6yT5EdhGVxyc1SPWvw5P3K4REdTiTdnyKEIM76UPW0TntyavTsaMIXUYQgAzXxF5
esYOLHojq2WDXMBugNiY8aXdGivN8aUDIOcgjzjk0I6f9aK/XNOD2Cj/185wNi5orBxOZmxA+FkT
DbkqrC4kbq9U95VL7RxDq2GgArQC12l2sPqVo52j6z52OZBbFWn44cox+9asIwDxg2yqDrbooynR
n3nSr/Dcd7EtaO36JgyY+Lx22t5BfDR8wDT7e9MAQ8YGo5T9Pt2+AgTpKaHqByEQP8m1oDgS5xR0
Yx6unDyaO0eR+fCGTU8xnyZFhFesBnx5kO+duHZTgZz/YxIii4agMU0syBjPQ+XNnVHVkLhk96qm
tQUUuObh9NGEC2ByY1bJ57w+qCqJqr2ZUJnTS1He+f8TW4ik9Sk108BcmNvT37p6QxSxPkCiCdOB
gbNCn7EtFlX1j/qpj0P/kLoEway6XuCtCUGcLABbApao5l8rxWMse9tArd0YmCRA0ofB/SEPIIcr
RzP06u3M/Wx4UkS+QEPwxwNHatN649AjLsvIhle0cwEPB3ACC7qJbQ5YEh347Mf5sY+J91ZUPMuu
iJM95t7gaoA7t3V6gEasmBHlR1J1Iu4uB+ntuE3DrBXAKLNAPRc2C7VQkUO6OJFoixiDB9S7I8xn
7DJKWgrsbrdV7Sul0e/LEck0M5U3dqA2WedK2mxXkGWQUQivYzH3/rxs1EU6t21u5VXJ43SwqsBx
pqb9qJqQiJ7JL4nRsalCr0n38TqdrcUl+G35xWnpiziD9P5VXdFc9whBtncAv7FMJ0Zz58wz6CV3
VHmSWr4pJ/tM1UH0wqAqrMro2kHRORITxGSZlVO8ze9/iekJoyECC1fFrjjF/4uATXCmxmPW2x4W
vnuY68pryBosyLg0wx/XrPlu08yEVcaPvlHB5WsTlIRc1EXHMxyF/quU+yNwzX69Z2ZNn3OontcK
Hpz2iCCSp0uCduadq9ySKa53rX/r4ypmS2DFtiJDd8lpC+SuGMOwrfOn/ZiMiXT/SB3pZcBt6KT0
AfSZd8z45vGHNJRUHttyFBjn3Q3Q1c3WUbv58mRfDoH8IEarToY7yh1rtD4JPvsFghUJn9I50w0h
oSC9URV7yFJZtDKS2RKkgBtEovap9hYpN1USAzzg7wwBedAZeKGBMXKksFDdOGtHr6OFnF3eqaBE
3CHD4ivIAoOTKyu/b+KVvVtBoC28/AjqqVASzX3Rs/WAMAJsYZSAixGw/8ap/hxCwzXfOD6Comme
9dLwQhfCr3jDvjy3+jKUHblRUIHSuFoJTgl6UjnQhxm9sWIsSP6fwAItxicAgd7NuOyHzZMJUx1r
5IA5Ky265cZYqGns3lpq62IG2vbRJgZE/v4ROXbf/Ke/OXQC6TQdt1YweXrZDB8pJUXZ9N27svCr
4vGMrqqW2DPmHEeNc3d17nE5hA8Y3NekN53xtblBTeX3bp4QAcaD+dwecSVvesr4pLEvxRQWCvqn
7CFiUu+K6RIpfrpguAjMxOsmPCU2SEqMwz+6kBQBq/YqltbHgUFmaw6KfOss3cOM6oqroLH8VMLl
c1wGhvN2pXiwcujmATA/1JUPqQ1AM0Fe7JNQHhP2b9kwvLdHXavtUSwY0Za7WA9PBbCKcm4e5RG0
cZiM1yQWBBdgUWm5CEytQWa/pfhLmrswWvWSNFgTrPHw/4tKLfyPIS/Z2EyISmgYBBZTB3Zjd8nh
nrsnrWNA7arZichcdiMHYT6sQi6SrQljZMIQiDta9UIAyg9ee/DHGBbYtMFt4DZ/F0IwD6CIiM84
v2hBHZcXFcfy7Jqi/h8LCkeRKRwXwabK/E1OwIqu75n/foUUN8kq/Wpekb6yubyWM+xLpgH8Qikw
euxkOWsNUpW8ZhHF68aRJ3cBhuAjspl3mHF4yJrSJ6OSSERPq7y894cFpZ6+qerstR1ZNAOO9Vwk
FBBDwCE0WIBj6L+ALL1PeaPK5YYdYFeAlzGjtUIg9Bp09D22kDV1RKFWZHArwY5B6xZdPRGnjelb
AoWsRaAwwuPXNVUmShOQSXzwsRaRqxNXzuuD7BsSw0U1dRPXUriuBfj8j/zWiW1IBVlM6aw5m9gT
6MYQO9AUrX1rFsvQMPIhFHvuNyxcDclFFt0ZBH2vnhNbymUPzXQ/LIJ1rQvS1Hc3b/r5LdhZqh4n
wPn0eYvHtKjaz78GqvgJBqOAH8ZAy2YsDj/Yi0RgjuoRvPeMhz/leZqapcroO9nyTCjQqb1+V67A
3oHsxMfh8BvMVo9vExcn0AJIyquY0BqjlpyMSnzL40dl6f82RO8XGucYBD42vCGoyUD35WgSvpW/
BeaBw/NLGOHQ5vZJaIAf6GAxNyoRqbYskqwqlij8aCIP7YXFO6PFYqj/S2e8yPpcTPmch8G/+NWo
0FCSKIqgy/7wdttvA8AAgHRBpa78LcS/aq+wJuFocCVjS+Q7Oba5kaphCnD8ZM2LH2O9/wMw7Sds
6lCCbv7u6vBodSlbwQyu75+tn9K5lqAx+iJWa8zj+SOGOPIlMbK/I6iAv/A6BL6jKKe4Ak4BOq/Z
zlQNSm+Tmn914tJhVYYiYBGYeAgGvuhtTh7nTSV6S/4NCemanwxGwkCPeQ507vFdTBXY4OTQPs3v
OQfqYAFdw9Q2gbeR/tomykRs67bSQVxPT7s2PkD9RXFTTo6TiKaXHhOI6IrqurGz6A10MGicSWYM
rqdwy2StCa5ptbJmkk9V0dAZcBzeP1tYXCPRP+/VqK9fpMybJ5p64BjIvMV4lYJaY3l/i78IZs7D
SZU5a0PwokV2pYL3KFI6RdUwrjYtn8oP56wjdjSA/Drnmq9QPqb+bBr8GvaP1mOcGzWUD+tA9ko8
NgLsZse8hNCrZ6Cm6m1+EsdZB3fvXs/lvJ32GdAg8SlZsm/RlVyx4pqzg459A+kPNFyKILDi0aoo
NFmjIxxFNsSfwjw8cav0eUrFTftqruDxIDqoyQo35VBZUObVMzy+WDsMlUw/tUMXbGRuEGclgp+N
6az86PW9daOP1MVHtjuEBsRaaBCK/lEQFVNEYcfSr8gGsvg4bgU97tIT6AkmUDd6mUKzIBKNp5Mq
cfydalF56tIGf25qnZu107ZYsVyLAW6oDpFtGNXKrROwcZL89i539D00C/Rvshe8Hu8jXsarwF9A
WIkFThrHxm2s0rbGlstWIbKxrX1wlGbrdwRuOlygimm2ffcyyoyPjGTWYZ3v4/BIaj/hHfoIxIgv
f7KbJVrdMTf1nKR62ZFiuxcMjdPFWZLpnYiMv6sBNLaByh/pvrn3D5eOwkhoaCi8/xXlU5MHO5S3
UC3IVjmNyU2QytHFiy5qWe27cFtawciV9dYXdESAnhl6bPcB3KoL3G1sNZabKVpYg5PLc2hwcob8
CTbHOFLStxJ55v3n7ol6tIiZZKJsj6XlQuyJWJ0c3Ye1trYKiRERxdLbdV34QaEGi4kSxwaSt+qd
SKLTphmyRS1YNf7YabjT31HctdEt0RcNKdAuBfIxs7n8Iu62D9m6C6Rbpt87XW3GSw1zVupaYE/n
t9/y1Byk7nbnsFnbAZ8m1Fso20luqHbdaIoOJofUqw9Ypodv0PmGiClG+WSvTFpJsGEjYBuMYk5s
v0v1lXtqvSSn9iQo1z9C7gjtpt1I4bT8MzoqmlIon1fSPs8gUu43RI8/S25H18SdcwtCrj9Tkpf4
fs0uZK+LzhpmnuBEAh7O5Dn/cvjYnJCRgKQhQBzlh0Co+tLv4OsOElyi67RDmsV469X0D+8+64sL
uRGMyR89ck2bxkqJ/PNosOSWM3IOFhUVHekNjF+0keZ+BQMzWjQeHb4qC/a3fIZYDAGgzIC55por
bc+o5WvkXKD9XDtDNAMa2yG9O6Lu4aRTfktaMBsZYlTPBK5gAJ0n7l68qgLINp7QmEmVy/mwXpJs
LaJGN9L8hgSIwtM7xhH5QhTl2IzSg7wFztZDEo9Y9WQoNS1heWTO9vvUC0n39q5qGX2FcK9Wp0fW
Zxz8UrToGh9BZZU+Bad/vqvTCGLeodnyhcMzWVmy3Acgv0p1ZYHcV4QS4NbUHczx1kn4Wp/vgHV8
MRm9YOU2NbUrGrVceFz/WFUdxwN9/CtlExW0HPg6Ti/CMmsrSkRSEjnjCUZ5ZiVwoC3PgWhNVFFC
Yj5AqZs5eJC3qqzQsv+Swu/l0RRYDebh7V7vF2zlrfqWJqGwt0juTX3Sl0T0WHT7xcSrwP0/VWT8
/f3Edhc5dFIqHImmA1AswFfu394NE7k0kzRi3zGEUFdIsVULoAPAmTdRxFfhcpb7aExS+nz/zmQP
gnsZGTz0i5WKQtCMGyyiQppxCVZ/sgKxz4acEASihjFysBWeKfPb3So4NGlj8jAhnO4/cJZk84ic
leQsTE6gmc27ev8xmEN0F7kRVEmNOpw16V7blg8x3+9GsEUHufzJltQT5CSgDLb3LYh4Ja9Dekvp
RPmKzwQT0ZI0/qXw2Fddpt7c5iAhZxHKeJBWqG++wdoDCSNybZj2iI3WHep9S4IHYjCBPABW9vov
9vrG7ccKReFZ0EEJrq8mqHnYAHjtfCDQuQLh1j1KSe0nj2SFhgHHfD5WlOJ7VeH8nPLhTFBSuCBQ
FhC/ABRbh/CK6xCBipz4uxCzpPENCTscHiueW5zie/7bCbYr9XEN7CLe7Jl/cPzi0mBJ8B9kJwSm
qV76m0BzNj0y/hYUDUIp/wfqZUbddP7P7zlzhqfOUD4fxHsKznSsrRHSJdEThNK97NkSHlLwE3nV
foSAMT0L7Luv9W60Fbd5hFH3JrEtWR2f65YaHJCWeOsA7+w15XjUZU41BAei6M3NsGsslt7vTbfr
Nq5sQQ+dC7EU5gnbGgn2JTZBMoRoIfLm7alPsldPGmp1wC0noTn65U3BJSALw6wDY6vCw4g3A/Ce
5o+9vffDDAe0adHg0l7HAudXViM/1eUVy5PWHRbxQd7zifjOWKKSOglYRQIBVBu6tbEUKRaJu4xM
aTSXIVDgzkSfLuLifHeNARFGddx8sI1sh51RluejvfDKw7xlPg28O7e72yfet2FirKZPu946fzyq
mu9JTRUlidKeoBR6okhPVegKwm5dQWyOQZlWqRMl+fR+1ranNdgKuDMkLsBepKHRuqy0fdZz3Vd6
/JhnnVhUxTJrv3nuZ1CUA204NtVMDY/ykxvdI5kDjLyRCpR1dCeBslyIofkcn/wIRSJZLwT6gITg
jvWgH2DoyL/eHfrx/tBVEZUStNxM7PLMarS/a66pDCEeNXGibGwIyyHu1OnRvBCuFcaYp/9zVAFx
nop5F7sNX0668eJzkiVj7CTYap77gAQbxs8hZDslv5vRvN7cK7DHqg2eebVFPIVLaK3hP8bTXYaI
4SwVeJt1EHef92Y9073MXlipV5W10+dINgc3XmSa5TFhwN/txG2JrgQapMyWvozf7sYOeG2nrIbh
knpsE+Kja1zAm2Ia2dhSmkDIeS8NFtINXbHABkhineXsg9HiaQI/oogEDjY6Y8jXcSUUHDTJ58kv
pKIEGs/tMOFaIO/yNhBOodhMDv6MD/wRwuMtjhkiEsA2GQtQvLIn/DzXw+YZsQR3LOiyNrGUoNmf
cik6KbFM2ro82CdBwvPATJxfKF7PFieAPEJUlRw/wf384sD1eY6ml+jbKeFnptKLijK54QVpQqmx
j46nS63r50gb3VHE4PkvkQOvqOSZCYfsafsld2YICEXcuMVh7SdJoCxdJndXMqQ5qmWbsn8uUFVs
GV52yXrU34OvopzO+F/CCfxys0WOB5MCWEGiKaFox+GYO6e5/pfG9sHL7wPowSEBPCIbvAdkUASy
6ly11MDDdI3QBppJXFWd8RCmNTeo+gtqtQiwV5yakid7nBZaIsdeogd2vpkwj+VFt9/vHl/NrjE/
zLovNBhLrP1nu8VeJiG6lTxvLK5Vjl8JHk6HZ14B9D1fbNkIeMWqm6C/UhNxjkQdvjXOCSc0vTGi
helxjGh6SoXAzhZ+eDEleL3ePSeVlv9ETGj7Y0tTcDWv2TonDsODftXQ8CmWlLYmSbZx01Mvf3ws
iAAU0idt4WfRRlNmIfliiBF+awwCT6/8vZZJz1e0/oG7yAAHjNTlgUOMiR1AgOKO30yc4rf1cTij
nfWIz1u1k7zd2R5MNfXfJmbhwojBye2hdgML26YhzLiWEP0TE9vN96f1gPkaUbFQ/lFosRs1MKGw
WG/1e6yg/mQKrPWvy3golVfdNOzqd5a4SrVs0bAQIqxqhirzXOPTV4HcNGIdJt2BrkJEAvz4qPvr
J6z1/v/pgyX69CAoa8zgSt318qkhhneRTnPXHmpPqyDOhA0Pl8QHRKF9FiJwftSUIGnwWMo7pQGu
t6Mn39RHWtqAkFGifykqMK5Ki3ctw9Il+ii+1++WXZB2QiXwxSNYZErvArn5lQn8CRXHYwmo7qil
lXq/g3/KePctfPsqKC019yYiGCWHJG3vzZRaIn5LpZdZqnG7uhbzdgHfvhosm+f+Tz/kM5sJcRD4
jFA17zEoTnc2T5QmFTTA+SUnzOb/PdDYafVBlBl0XhmKFFgMkCSo+pu61bVO+jfxxuXRSt0K0cmF
oWj+B9qJ2mktVQ8N9oJXcH7+9NZbMnXcYJMa+3gDRhLCpzNbT/ONfrhLoL6vAhssMJ3rJU5wLpVT
+4TFR0pYHtjkDSLVuyFaGPcff7BY/0nXIwiPGrkdZeQN+Mh5tnJhW2xcxrklWOX9kiXKh0iFRUDH
PXNtQNyxrBi75y/gknxgXu0t5sfKwcus+bfcwPoMcZIq6h27LnSw/WBYPrzIOVOIYpdLvt86ey/5
rUzjr6CgO9gwmeHMcU764wOHmdr7j0i4V6mfrJsOQ9vxhDhXHJtZ+ybAZpyI78ojgYW3lxLMlsr9
kNG00czllSqgbcA6+4bGqpSOY2+D3r15xt3Y5EYLn4ALs/Sylpyb23i4pzreSWyXzsId8QD5g9FI
A0W1acfJ/ieYiEeAPOVKE3xy4p4mIZYWU51hfGzenbKTUCMjimlfYgvDSggasEs+6c7K8M/Ed7Z5
vCNVNhnt86v1KV52ajZ25yW4vVLKcbDfvqTsFxqYmoT/nu+23FzNlrQU3eQzH23zaqmCy04+GS0G
EWsDbge2RdRfa+PvqSOWWVWSQSMmuTRzic8pnONkVJNfOBvgQqeKHKJkSq4uCXP7Svi2AzF8c4ok
R0PULT/thtObI4hSJxqOwzw2L7ra9klAI9bFe7hrHRjOg6IfcUzn7vtJV9tBcyA0hkv2x2SdAh9y
qqOJzy/GZMUxIoP3t5EgU5SlhgJvw0nXpcUUJEnG34M2I6qjZnYb5dsYTzFekQIGJTQT3PBRIlo/
y9/QPjBl9uYnFkn5hO3EjkObJH9ChV5CzcFpDpG8xenCCSBby8DuDk/0XIxL9NllOM1Jbqm3Mtbh
L7w+oct32vbm+qk/rRfVh/PZnHG14DnVt7BhANCOKl1plfWNfFCWZqAbfMm0oc7gwBBlQpv9icr3
Fel//KXDxb5ihrLfB7rKWXXury1hCKE8gpCOoh/07ZlxjeVviN6rsA5H3PKWLvp7q2IbDYUkImcb
AvuJCR10KhIEysn2eIGfeA8AEG/rPCkrrLHHbSfWbFZMdnVtNtxgFkspsIyCCSrkc7lvaRoQbsGL
AKW6qL4/nYsMX67xM2sMQooUE4HorsrTnTPIPaV+sghN/yB/YXjQgG2L8dpwKOKi1YSUXpmVf9oX
+PHi+GucWsj7EldmmCSLfNNUFbMsMrGjb04vtHSJWFbZ3tF3w7H0zSJOQ9lKrqbCdVf+Q2TRgD/4
XI22SF06BMN0BXtGtuXgl7zJRjbLhXVA4dQyQ9HMOLzNAsBb9CQz6xnpko7+tffKtkob9emFj12C
UTp0QXqS/v+1/osQ/hu455gJxexd6ipQF2KITRATMwgQgmQIpHf0yLSBQR28aorfF6f2kCIpF9Ve
EVQjiLO+BUup5TweRNdoLcfnpKIBwkbvoOQzhWzTC72HkWqp+HtkNuWVvYMN9yc57qZ3A2v08waq
G+PZ4AzVPV391We07UXCH3GKaOTk8x41BNzQntL4962UFuYSEq2RbkXB9aF2d/ACYS4aGqDykE9g
dXqeFoZ5uTJd7y9TW8wIBza+Hs6VtABptO+muKe0Ym5NMubx8Sp+zDSDgv/uY3y/ER4582e6dknV
x1QkSnBTKbev09YH8DjRYH7hGl6wSDOwznPtUiSrqcA6npCGS2qmYUf9HHkq1whpIdEy+U6B3cTA
N6djdrw8rJfOATB+wZf3xX82cio9l/GFxflX/oAaF7uGJXKrPa03+464zJyNAwcr27ZOFuXjun/F
OBitZQirNvxgFRn45JqOh5JSLwbgRAkeLF8Y9R99XJ6lE7NbGZsE8QmnKnuQmw4Ue+ezCMDC998j
1f8KvI6g7oE570kduv4V5a//WxRfWlHvfNgFw0SFz5mmUcY7WGd+waUK+1bRMyYPucVk6jbZYSSi
nsDvqHtdkq6STQpEBZEl8BCvG0jd5cJgnGG52UHKKhjV7HUZGCEAKwFUNj5Ybh+uu9Yq+YdSSsnt
iqu6y6WeRJmXGKD7fadgOQbb+h2ype34hDzvQ7z5YVZMgpBaE3XDax8sAtnNPlhs8KI/Q80hw59h
lqzOvFF6Df2+gcE5IpYKC+HYtkaSYbRJRoQ5qLpz4SzbUYs3XOcReMKCz30OrpbifvJmTSTc6Jlf
hxZ1eSmUelejt+tlhbaFcQUBNWhDDBMHsl9G5TDwZoD0KqiUA87sJ97ccrIiPQ80ktHhhVfIrGmg
dUVS5k+wmi3xzE1M5tt6yiYv0uleuyGFfYMbG8vN6iYs+aM5bcdlPiS0KPA9kRurJfiNe1PWY7eb
/znjWVY4107F6m6HPASeZjS4pRYeyoCqWPdspyMYtMip8W7UjD0N6L8WzvJJUg0jOG3fA9taUyZb
FTJfcchbOPhhJjlqmkafIqVQpQKgdehkOX/olggoEqVxOhDhNIsxgbhVWMiHxTNS6p22+T2voiKh
93P6/Rb5brx55QpArm9j6vQBQ7Tj+B2esTKeV35MbKHCzWAFsPBvTo90vsVrpDRXJslvOmceYbyN
fE+ABeRA0SRX2wo3FBIR7jNSClC/r5hHt3tKswWMdfBVfr2KZdabZRIuTPdJshVQbC+rWXfLyI8s
7XWTnNS5LO0HtTibkuvhghpLpj+o4mkS+U1PE/lGaFmRah86hGyfZ1a4COdDELFBUzFJ8eedeJPR
LLITqm1LmVWJSZbbjSz9FBGy5IYSub3Dc2k/lcxxYbNnR0KSPF1Fvaw3lnLnArqaC2r6pnLL5w/Y
D+o8vL0h25JeC+cJe6QrjTY2Wc6NV4TQaoCaVFj6BUf0vwENzlSwLwh2VMMWM1qaKv88411RTSbQ
1ZFJx0UpSa1X4mN4UqoZcH+0/9Ix9X5EJG7X2sMAIGalfR24cOKWzLItdlRCrHCSFwIcVGbfnn2O
XL2kBv/OUq1EHXn1arPUldpkccRwrOQZcbtxLCKNHb62rtNwCe+GljvtTKo5MnrLx/d38VfF6c9l
nwqrBBA5wcxzUOXaJIJ6RYXsBZ98AmgMyg7QsYIpNzRgihpH2k9D27PMbmg6+TEROBxDw3yk54eB
c4bfebv1sVH/1xjF7YXtrLcBv3e7KIWr8/p/VJN1RrBaXLqQI45SLrUtfIOjYT9eSofBqwIC6d5M
dIpcgY56svtLK3+Bm7oYrsITZyauqaKBDVeaKRTjGfBmdeLuz1u/417sWlPXn3PP90cGH0+3iMRk
pEafOJD6SddV4zDZsIdc0lOzi4Y2UvvFNv29453HRCwfaIYoLKzIDPx/vUcFCrs1nnkqW8hkP50v
hq3h5wWhBtLNlVn6uxFYhz4IwaY6pQ8VUPTdM7coyZ+ucDiHd65324lpNg3FRmuTkH//T6ptCvkK
wNM8tUYFJ/HJ9iLcEnfKakhVbXRKp5pZg5FZRCTpQJW4eBy+Dq2VrURGW79KFxn3V6ITMm2LPlzg
CK/ki+OTl6oNj/2FZbiVpKjdhOyGeBrCDCsUaLMrylM1yQHRa6JQj+1KLy7u+LlikB9fMqm2fGUH
2bD193J4z3nhaakP4kyjbqePDNXrKBXFZEOeemAn702qf+Gg1wYECTOLsGnPVmcxC4LFaiH+UyBL
Fy9UGuEDD1D3GqfpwHJMyRw4tJAZ4il5YB5KzApyPcknW9zf8C70eKf/PgcUf+0djM1ijnSG25fk
6E0v9t0NttR+Brzm12nOH+6X/RyDjUh7gDdxfR/P2B+wp3PY49tlPfvZLY5uPAQBja67jX+Y/uFB
8S8gYQjKQ2SYOk0XJXqWzfQZna8uK52hsJXlEFNRaHA2h6zKVGnl+ZIFDzWoO2i6bbgZJQcPVG6x
wBLykET9Ct95YChK6fTu+uxScGupSl9B+F6DwvR1LLuygTca/KfQyXxe/zv2hMBw1tYvrwq815ES
67lVWERbqAMF25jy3KG1knArgFQYuajGpraRfeTLuN9BX+KqY4Iy0WMgGJVp71hndGaaN6b4u1mB
3gKEGhFeD7Afn/YZLVUL4fJS3RXZQBKgvEWd3HhEYe+ZMD7xmUSqryQ3cV5Ii9qGzzNM4aZ8SWF1
2lb4rt7f0KYxDMOKyMzf2uyhRIjuQhuCPuMYn6mpp8NVCLCvva6FnwostD92I4Nv2SGPcD2NwFfD
ddDsV/pqlQOHOmhB1U/f1sId9Lrh2EsVO44as4OxvfaXrIiaMCBTuitzecIaSLWvTG2H5B0HtUcL
r6Yq71j330+pfbWdzQHHjfHDLGK432T4jbz2iXbHOLiw/TeKh1Vgg8A5nyszwiz8QMBnU3+VdzC4
USjHJDAg7W37V4cNeKPebiIZQYh4dQ2rgsIwKHiLqrStQKZD2sJ4QtzCTllASc7WuUT25xdoLW1F
7xPCbydsHbBmKcETBUt8L4+8uUbh5t8vcZvCPpDbJAmrnxmDU7lPGvdd5Tpehejw+muE3SGifuEM
8AHrkaQRBY/wPG7LTQCXZgtvsRKL8OqdrqRBtNBW6zbKBvvd6N2RB8VU3JYkNalbs74EsFGsqtEM
+z7XA2spK/m9fCtJGJR5Go/AX3LVeYiW/Wy8PRuQ7eDW2V73QUJjZPmMTBUMBeHeP2Zb/aFysii4
poZ9+2PFBCgTV/lS27YHa95Q43Uh5AT/RkagWxgq6iCWs962jUl0K5OF6SYRqs2zGuCrdzi4W2p6
YNifcBnX0V7MWKhZ6hM1yqfZ7kPGB0yXnMG49vE/aMyU+LJ+nNUPcPzZQ5Gl7BMfKxNzsihzouUI
TyHF3+Rd0DcQisDPDZWoOXqcXPnOrd54pUGVz8ZZ0A532nhxNuwMvQ8rB4/fQwufNHOZGK0tEOsh
pjLrYBLnGEomMoBZr7Q+VEq+wwnbhjGA96j3CzppzYAuqjT99zjz/pYzxSo1OBUobLXR0WK6laSH
aAN8eRloVeQnOZ+JeAMH24rTGyFJc9UhQwzhQN/gzA1HGM+SEx37H+F/jfBsOPmwdNdWBASB98QJ
+ScEtSjGI+7fMt65Rlf1ZJIV1VulMZzmxt7XkVnrrxBl0v1iwzKSI9Jo1qryEXPQYF3W9qRlApOn
e4JAiyCqBBwhZdx9U8i5c8Gf8pA9bUILemrzprxB5qzn48PJxeV54UseABLZEft+XlNT5lzHI7Bs
GKekCBh1KydriIteFCauxl6vBzw+2WBDKMEWa7B6yhDrUcQ+fcH+BAKhE1Y3U27rPhC9tzzGIx0M
MHzTpsGoBcRTwnMKb53V3JZBUzuRmy9SW9jU5WsFtp1bwQ7IYNin1mCpXEz6zYjerO9lOVk/SEin
3yvdg1ynJmgkU1p3YQbh/o3+nTnlsv1FFbAIngdsmTS13tMLeSQAJiN6a0G4naL+2RjSIetDbtGN
DA/XWJudj2sCPj0cSH49sAz22wfdroBe0vJIHDla8hyt2othXPjSAAzoFpcc2EkNI8wh62+ZHF+b
sKC+phj3ajjhbZ7+fY0RXJD62p5cj2D+lbjJhqYsG/jNZEwPvIqOA6PH3k7bGSeLVx3vHzbxEVY/
d6AtroIKN4S6mZLWKpfXmg642A7JQ9nXvjfVTt0zIs+m9IdqwRHS83cSmJAFBeTbLOsrd5X6a6pX
/Ia5/cM1qAJ6gwaf4qxnOKf/nlDINz9eUsMi1+8KIat0D8LdfNt6cSx//xcYErJDEWxO2iTVGcr8
c6OY4ltPh9Tq70ZijzlamJHqJjIJB1lTD/pCrhgsFU8vxkppqHmDz7Me7XX5ayElt+kvAnkRbiqS
EJ+AIDv9c5AOXhm05BtdKt/+9rWCkKdzLDecSUS17qKWd7Yt2JFlboq+ndyj+P7f3L/FD6VoPkyR
yBqnGkcDa3mzZmEtKjkzI1dMFK5nJWCFvV9X/M2hEKxum72F4tAszd1j3gLS2FZ5+PMCPMYIFThE
EPmZEAake5od2VaoaaRV7RF/DCKYrF9Lt+/tKmrXsLKEqCqOdYSquqK0FHSxW3E38ET0qUyyHAyS
SwTNzZFfGWUPg1j6R0IK98z/eam9DiJPnnihP+x9/NPJc4xmmqsMsNru0O6WqHmCWdmoM+8G9zNa
4ul3GFNpH8em6SyZw34EhNg4T3zBYUBtZvNbnGsbPIexkQPT58D8gfDqj2Kiq9bAG4r/l9WBF3FO
LzqHRwcfSUdd/mtr4amRwHnTqhr6W1bK6GZt3EhaL80O7/CNQ4Ukx5ZUp20DtG2fAQ5AHXQI+FnQ
MV+FXuKjgHxuT3QKwg/ZTOnrRJzW+x9rp9N/n5NDdnY8o7R7ZibfJJLXc9Cg9HYd2Uo4LznN4m3/
3mMsSPBJOWbq4V3OvlqV33Vij7eqjM9vGRWZ9OHnkqSQhKj4cOlqsEDI6568i9hjwZIxig/2H+Uw
2tlre4BD2j05S/KKMRhy3f71Ha+AWmTQwFXQIiYJ0LJGVmPLFlyj/cJ6ASZcWX9jBvBUYshV5GhW
ymIReNHqFkF4YCMhCpRSyPT7YmSZ8koo3M2LRsL3hCxrpya+Y+5sCk+rrxPaog/3DBWCmU5mVr7Y
UZ+ylzMcIjp1wyZQVwbq9+F8QPBFl9t+QKmi7p9WxFEUbM0kZ3EaPG+D1YtV5OuHN38j8l4pDkuf
N7TKyiGJW6LxcL275AhC75bUQnYXjhp9HSYjzobvxPnOIPVkPxUhnjiUo0iM9BoedMxyeJUeAHf9
3hlvp4F94gWj9/opjBkulVrZ9GnaanTUYKHcPLVfejYap2p/H0ZPNnwDsr533h7dO3Sy1C6tP8Xk
Rw2eWEfA1XFgec+EEtq4NVTEeN0mPxfqWG+XnLlZaXm+6IBhxniwYGI/6DYjCsp8OnCJIugpW0w5
fjUMQk3udY6D6OGCZPqg710voOM/QufJVD1+CKgDNs8UYMLMIyisvEEs3TyWpDkdWhGxcM+iPx2z
aqzLzkg7VsnKsrrOIIqjOG0x34Z7piye7ENMaFiArje8psEcWWkfnzkmvrZ7L1JksGgqpJslhd+O
0iH2YriTvK37e4KaQE+kYWeuVN6wpxhoWRTvEVf3+41uD8GbVmSTzxMH1FysJqptzPadosogiEcH
eEUfd40IpplA92N6QznkE1CxM6D2qX2nRJIrZ9aL9xUp0/PWW+niHIZxiUhxxKiYtcFRmOGFNLaS
50j4Tz7wFGIdiNCOIzTZREJEtKdjm7fbNZbk8rAsPUirbtfxVqVmQt0dIKVVJ/AbDMGmxbV34QSU
oKVgZAUsGdf5zz4HIwSRZhSuzS01Cq3iVqX4aI4g4o3xjSA8yq3BmTfgxoX62OTD0e4nHZWnBdIs
9xwE7Ucrda9wLh8eqTRwaQ/4Ty+hDrEaTO9w6HSbxODIxls2QJy5SnBYWsiG+NxY6dB+ZRfbVmMX
YXq89k+nRULhdkmJyRp3YkUV8uiaIgWlAcT/9o/JYIgXw60wvVW0HKqpAWHPzFBdL2nyuI5LsN/X
GaOhgM1zQx+0NCtdqqQRm6v6xzsN3OFh8CGw4bawNetkZpaEV0laqzmOXUu6BSTWaSa4TnobdrSw
S049jchGDy1raGkH+sjx71wvikAfZ6jKQf64D3g3VSkyXitC4SeDRfQNlG5sHatJWOa1/ZHJK1M9
NFpP0HVNK4JRZnev8M+Ixt3GJNru8gFcVkFd4jhUgj7ltdv39fDsWhC/4vkNXgwh3qvwMj22+T+4
61JWi5Ya0oCfKoGOCmQNocgw72oDaRBxRJvOWCjknBZ63P+xvWJdwv3RtyybFHD7azOXggPrcmGg
YZAdz91lZ1cRiJqX3rs/KtLr2tlL9K116/wOzABBh8sISgNoZTn7gGlSJh034zh0PIsDT8GKHleI
Ehc/+7twg/ZEPA/GKskcEyDZFsSnb1zBTwwzHT5vCSbC1hw/sbzaMAY7U72ZYzy/7gdY9XoBaeYO
NK9vfQjii1BnNcsRNhrdW6UuMmhb41hT6wT2wit+o5InKpcQsDyfrPvsf+SuAbLEmy3dsL8Q5HUT
nKtTaQgH8H0jjO5PlzoKDueZ524m6vviW4Czk9YPJi70wNQvjY3bIRLT+iIrusO9yfdT/XVfs8C6
YOMTbHIbS0EEifvVALLP947BjoICG7cdXGJtK+ZkpIIZVhdJc244bAh4mhzA4l9IPMJXcTnPqG1v
QbOljef3e2ssmYGPoDBoZ1iXInenaSMnUGCoRJFkbg/JABv0QQ2grmnDo0Bm4T2iiIXT1iwWEoYH
JWxM3vZDY3qnvefMwyuBJLKKEKECK2vH3x/BsDM0Zjpfb3LXj3pEiUiHtd0Db+HrgD5wrbw8OC+F
s9LdImnuslIwwSONMI2Yv5ZwsvFtz1v9mTGkpU9/TYiZEAPdY/9H0p37sMz8cEKvUXFHl5GwnB8C
BEcQaTqkGut6RbRb6lpjZafyUfhr7/TXREu9s+pyCox9U7AsLhgSbwGjmisl/+Asuv61Aihj6W2X
rpFvyywVYFnzNTFHN6ndt21Qxl+5oYn5+XysWpktNNnmhlELm2R8T5hKJE+xDAvfryuxLmaiCxMJ
u+c8vNXBFaue+KVk5qehE3Q1WDWjS8l4wuCuXSUOiNJvpfWaYuLgw3odUF+peHWw1XepPN4pTgzH
N+kUAiUJQyWQXQF807KJGDMC2kDHRnWR7G4YIMPL48ktZdmlOf0l6xovyPwD6258dfkHSwtXYJB5
cBXDB/qMieiT++K8Nd4kzBJuRkAFmntgrPAAyCpLy0ge6ZZK2on1lzxN1SmtfKC6H27eGGxkCMuC
Aj9zEFHCnPgj4wY6tzyhmOK+M7b3GdkQODNG/txd55CMHpKvOw4+puR9JU3lasDj4tdUuXTmAgOG
YClQisclvbpTQaDdkmxh4r6O9b6feYeDncusUE1T8Pb4Bz7MbveaR23Ff4eSENi5g1hPW9kg452S
YHnBTecMQAnJfggTq6ZOem/SZ4NeEBL9yrD89im9RZ/cwt2zHLI4T6gb6TZfcBrNhkG45iBF+nxK
nLDJWqHGSHxQlCzu2YNB8GH093z61jzu9ACirosGatlBP1PxgXwS+ibO92mx/VHKh96xWudpKv1C
l0WApgm5q2PhtbEuWKtOL/lrRkDknjf2OZunBcAGy+Qgy/tJ5QNfZTaoXj/DwLZdT66OSiig3syq
yobyG9R9bMOb2zWQs2oLerXpa91z9fHrkIjHoU+SbzpCYbAZ2Uns58sS5ltlwNGCKSsW9+EgOND/
dMDvoJA8U21kuKMfm20hC9iyiXVWTg7XzIILpeYlZJ1agex3vOTdSXjSAMazCAJP2K5OXfNFjrg2
FPYsnsGNc6Thcd/1DcZOA7uKraUISV01Y0EfN88vzY6KnL3+6fTqHeGeUIJYog8yeBLJzrS8j09X
SwRivSPe0cjv/KHP0dkWnuKUcMGdGxZHSTiFf0tHBJMxvQ/6AJbEfOu60go6MDdq78RZ8WUDe1oW
d7x3bsZ8uXYLO9UNkSlSSRHriid0jK9QuwXRqcZ0ACIX8ibQKci5ZT5pBefanoZKCeD39Fwxbnfp
6BUyNxlc0SQJWtDYqBufT8fJ+HT5+DHgM5fPhX+PKHXYsovjSUiDOAJH/OUIvT8acPWSVp8QrNLb
KPyYBr14vTXMPCtsPYQ43eU7sEozGsowMdBikvxItzrOumjpSPpWGftIeF9OMfRVxB+L7RVcbPJ/
/ebk6AocavnvRNYkZmLpQoA46dpIxcWTv4ho8e8J5XfZ6Oo+Fcr188oVLuOB3N6aqbwHop+eGULE
hE8HUVKtGjmnQac52iK6jxIjIddixb1B9wtdDT9ti8UC9wR+jKx7LzWA7lA4mnxexsBsA72N8iMk
phMvWk2TIHaBDpRpUIxPQlZhGvwwcYXhWqlXffx4+0lSkBj1RXM+O/437LU4CGQN6h4dftXQx4wr
4noXP9770104BkuRPvYA8KiSML0ChpPuSFPYQ0kL8hPVwUCtItjVulzNy5I590x4BMfkcK3ZFbgn
uHSTIvRkhcOBIQSe1SHfouB/ophmYJbrlxeQ1DNU8LFzhBSo7tcLKMnPKV6zx5WpkH7uEXs0RpAy
VCTwoX0O53J8Iuo/G4v0i4SeU071lsYECoAll6gN+3gT4ARBFewwiOOAuQ/c+5U+FEPG5jTSye7M
4TlKGihPbC70DLF5BGJZZ02fGqNc+tc+ZCWQC+27aBSi5Ah/xkefnGa1IDFxid41sF6tSfGXe07i
bImHORkx7aFA3+TpNKDPNTnabx3jhMMYcwC1fhWMK5p2n4otGxbS22dbf0awPnDVD1mQvn/VwNYV
pT4HS23yo/zbP6s08PHRaYpuLJB99WlHHTCNokLkIgkWK/LLAVQpfyVk0b8B+kcm5ydQ0zxDeG2n
RK5dDLkiWxWqL9GWsXlnMWZYRkZiAZ4IdcqAZzgJbHoFit2jTKYvXILboiOtcfO0AaRMU8wjRnsm
yZj2LgfqCDjlyGHQ1soxF3Guvum/DOAl2BO9YVXP1LDwPf2jLDBQfatUlMoozmUdzekXBw2/AljL
HDmDxRpS6DRGZQR6oyFfXz/zEENzDkiFK0uC4vet3G5wi3rgKal8LgYcPdkHBm/pjxFcezbHHgHf
JRS5775nfCfBDiJREVKTmI5pyBHa/b5n4SQ6chdfWq1M6JOm+7jrm7LIZzmU+YKATTd5cYLx7BCq
aKw0fs0hfV3yG2C/Dm/2H+cvLFO6gBrW4+I0xWdBr80PbPYGrT4cjCFz2FDN4g0v7hp+/HAnxa8j
VxjXNLTEbFt6xTySZ3cLV+wV60Wt8ErS1bUPfGQoejdffMoMZ43Pcm1Hmd9byY3MwSEPM5Ky1tWr
7e/npFwa1SG5nORG5qORx2PAYOgZi8N9ydogvSTGc6I9bttXqx7JFYeX9cUqVuj3sJj6XzIsgWja
n7VZcTrGgfnAuF91xUWnLpEj6/uP7idY11b/4ZhsxgIdgZ8h2rH6eoiAM/XDL4alpY5wyKcPCJFC
+2c/fwWNl7WFY/6VOvODiF8NETb/2upRNQRoL9GlSgaUAltZsB/P8yZ/zTsfYFM5d2p8KsRmYB7R
XG49sAfTnI/6KbIkfOwwqVKTGirz1IGbmq/ZcWE7aawyldnY3oa0oguAKCScxwOfsgjFzJ+4+Ftb
m0ka+RWUP1SkU2XtFv+YXjt0V4U30aZcuk3K8jKsXlCJR1xDot6DjsIkk3YRzFfwzcgHkT+LYpDD
JjMcVgXDmwCXtBnK9e51O250L/qd9tnnnIbGQakcV5ZnwcS3yqFsEt25hJNOLovJpI1UBrG43Jgl
XvWFnFRmoBOtQZC54XqYGFkAQEvEPFP3Fha0NG42YBwar1XTHL07n18GPVNdiSxQZ8IVYZ3fhobS
R98ARmp+ZuKwgQfNHCRk2hwTQQfBBNlNzAWGdC0X1UyyCYGcn6TGcEZbLrSIofoCy6oXxG/bHMnC
Bm5/Okyonzx6i8A5j/Na/HcPzrvUH5evSdOF0/nUS+3eFlfFc5Or1MCBNWJpnDgZIV32VXb8vHvj
dDCCnkVWgYN5NrOqmGBvW28f0oDkONFcqPrw4IaWTEBxh0I81/+No2c0zOatmKPxqNVN2LWu+rfd
9wk/C7AJDF/BSr0YveVuP7qA27DSnA12cieJUVhs0JJiJ95yLKRuUVpKwKc+UB3s+HoK2dloZ5aL
GdMxWbrNfAwUMDPWCS0KwniBmSu/D+w2i/wGuPkWyOPvPtiF/Hkg2DnQTW+9IeFE2pG27dGuX7M4
JuruyD5U9MggUkRcNehOJ93TuwsA026I0qHPL0bmWCEtMba5+wswwL3aiUkKXlEpOG3/cfZ98yX3
4DWpsb9oxzzqFnFEWdOjHcWRa9IwhNKNy4TonTKa3W3HRCq3GlyKb+fFvBPZCNxHc4wozEP/TW2I
ZPficAZaOreUlX5gxrhTLZBT4KQK23huTMPAEv6FkyOruuenVuWMmTozYfYLGVvX+3TomnWE4Yz+
IQSGtUo+aOGa/6DWlgHHtFOsUwNP22VmRL9EnFPHLcU6KCywLgb0b6H/+tXDpvOuncZPf+BPzTHk
KPC8Fdg0e8tnIpjkx0XkAHIP/kdxCykInkU407rNje1ZNFGiScL3RIK0Qu/48AOWbmBpqqHUjZQU
RMhT37StI451H3j31O4RTk53aa7RexwtvpSWEj3/VmPIOly9TSc1RxohgLIrrb7KagZJaJYPPiNs
jol0ZLN+AiPlIijy9lfeq6fhiY5bcH9NPOuPlKj8IgqU8PECbYLKQ6EUOEFTWpJxooc960RyhXW3
kRwdFmcQ2aezYM0x9iDMi4gcMbhwsUYnTzrKqx++6RJDGEEa4J35Bka0bTDs5AZDaadvmSVtZOuv
ZDUdzXFnCGH7NejjPZjZtg64MQ/xhgQRUxlygSpNn8I4BOdVGAINNEb19tqKxHYYiPh7yYKYnCws
6d6s98hEbsp6qMK3J0++tK6c6XaaZpT+gXINf2kUIHxf0QHSrK0Hk0NxwI4uAw8h8JBru1Tojuhg
Jkek++hSfWOjMdm/xByhl4Oz8voXHehyHWeq6+aJV6pA5pBP9pbscsllB+uEZpDxfpLbYHXj7jVe
WiRlv/VKCoSADYFspmADb22qTcPVqbF9XfdtH3f1vQcLYf7Sc++drmbFt4KjNNhKmhTeeJit/E/a
AYpSANaQXh88hrhGa/EMBbt1mED5tUwwMdUmyDiXFStfjDD2lsdBg66/Am40HGOs05WaQfkiJt6R
9IKP/Ekl/mbZg/X5mLxJUpWRj32+zzpn3pZTHaE79sTyKUI6hbcmDWQtxP9UB+jHi7/YPnlHzcx5
FCyt5BWcElrgqCYitKtK0msRdOqQnXhqw7SHMvWy0eT9bZH4gHtvIgZq9YxnE1HoB23k1Fg62hkn
U9bPSX+/ZaNat3bcX4nlwszmcLv9T+s9WkMlDb2lFN0WpvqashmDYsh4UlJ5hUNQjIk0HuT4Mnz0
siLRtC0mghmZ5tV19zEvRsQQUvRVQQmuDutRyC5Ozqh8SVXKMJUSrcSdtD9WB/1H0br4GfgbKqDy
itz/R7JQCRvQr/FcNp4kOfGvB83DrvaKrRQeKMcScdjNMesXQ5Jsqtlaw/AdSU5D4wDrWvFVu3TC
TkMb/GQnPA94I1rZ8jm6c1SIVINL6tsXI8Zbf4KnccpjAPKXzVTY1SglD4pHw/DKxSyoNwgspTVF
SqkFwvyYxwx3Zu+5V04SQHtjjA0sIuLYqZp1NTqRcnRtnEU72qQ+LutwU7zuv4AAbW9dJAso6KyP
Jn3bh7Kh7m2Ng7ldZjsIIUPPq64FGyt3pxPDtNMhcyeLfqKsFNjWcZswYl8qZto0TK9tCELkwmTs
rWmdWOD4w2xPGoeQ0MiCOycTMyzdbwCNuR5o0hJN7/JJIKj0FZvUcVdNm4mIJlYknbrrX15cbWVa
ESgEJ5qfBNdi0CgBzVaQsrFtd+r0Bp5mxODBGDuVIsQ1AX7AiDJx/E0kmacV4fVKzxmfFPPyBAak
rJLFk5DbhulnwOQUjEA8O9639L8dTCp6NXyfa71xPK81zq1C7eRyFRRPa53yiyXYgQi7yT9bL+NV
Cav7NTgvr5cDqjkfsp+7eU5kQfTEitRnK1j/KM4I3OBPIGURhV1M4hQCLUWSMlxbfQYzLsP8k5Ok
5y2QG8HIfB9NtRMQgPnq6oRz8y6YghUy4bDehfu1arWcF1v7VFlJBCeErBbaMW3po7oSMp9Q4kGI
+sXN4L3od7GITI7DfI6a5azPibHtgyx6tsiTsOaimgjTKG+BwjATskU8EAlrvUoj4jhPeeHK9w9V
Dmemt/a5Z1dN/qSlu0vAQq8b/N8DRJ6MfATRXzRgw0J370nGKAATkrME9jFb/qiuPjSNcTtu8Wmw
HogLrelaXa4pmOJMtgqHX8A9CEpIhFppDFeZqyfQKyNzZBYKGOTdrFD18HgoPG7lBoYIa2US5kA+
s+AM7m0hnIiI2nMwxGLPvuC67tZY1R/hTFkRU09gqWCGociJCgg8pUAGyipQEbIDz6wox/MtSp5U
yaP6wFhTiSJ8AxRCgzyo287e5RgmCElq5/V94oOwtjlrH/FIbH47wP4r5acrV4bT/rE45OiIOqRU
C9rPCUi4YypEFYk+moNZFvglQ/9P9ogcGoK1TFIjwvtgqwKIQ4sOy2FaQ42wASKU6aqj50RF8r2r
bLMtIHMPiwpyi/dHItpzw6paJDZAJB1LQQNxoOZSCYXbQ3WzHYsPUun5maMJDtA49BrlNKtPD828
pPHLuNG2/2ekLwIN0GzK/olD+HJBlieyG5yL6gwmU4OOYYdd7v3kJ3RqSRE7D/QWS6QowPUjQwhW
qFI984xaHh/webKCl0OTUyrAcaivsUMl6I9t1fOpETzGdAQCliN/G2GFLelnywagW/YDqKr5sW+R
Hpp0vXTDsf8LO4AjP4QuG+UkbREv3ir04PsjLXV5/DDip6dGCu/4PJb+N5UXAgtPfRfI5hfiMesc
mwv5+T8Pcyg1mvRFHjF3NaDN7lw4aBPDEGcTgmJ+XFssi42C0svppjzH1U5XzUbr3Kt6hLyoLdZV
EWr6V4KlUCRzcpAd1vzzq7rDwnHav22dU1VtrH2Fkw2l4REs2JWIvKICPDI3wmWa7vNdNbOwvbNt
jpsPqFkiCBbOWO8R/1PZumLH5C+kM4hZT4UVCiFFNA5dn7MPxCrH18SmdzHbmx5lHo43SG/cXPPD
VR/BfiUxGQEAMUZQ0/hoSwtIlu0qLvKYUoV20dn7vGkLm3tNBdbcFk94n0EERTfOdWPS16vYtJ/8
X3s9R0en6JHOEtNawae3UiZ1wHRu6+xYwZ7XLoEMNvzNJs9J6n1YdgQpoGZZ31EgF8JfwTvVATOy
+ZV5hCyUBdliS/UWJ+j2Mf6rNHazR1H3UnjGVP7ZYa/msUW1UUjksAyXn2FdXgXuNXTYZdvlCuKO
fbUqZDprw4jtM5ulcGXdZpYIFoA5pK/6lDLKsH5cLeeK7Itn7FaYFK+9w9wS2KPYwOYq/I6m5UBp
OkpG0G7U3injZnVkqtx/MBXPP/uGpkDEDHQzCUm3LVc9o79shEakJndYNFrOu0BrKT021hBDBf+k
6JnBCv1DTBpRGTd2mNV7AYcEYZMpLcL3gSKZFVz9QfCfpWwDWUsw06mPxCCsraSuHiC2QToBg59g
g+UUAnClJL5bLiSrkXwm0Fz2ktI8/6rxTbhlR11PwAZVoPunmfe7A7Osru8UgL8pLZTAxpqd7tpZ
OBSbJn9UQxRx1AXyO/MmvmcU8Tcb+Rx8tfWYpUiInrZ9v5sDDflRb6YvUVro/DvAyElx+jDbQk5U
eaTewV5XLUJ9/dMjLI3IIR/h6+WvLPsotRQLCoTg/KYyD8X83jgAyYZAeJeTZ/y9UcHadrOJTqD4
VttJVP/sRzLv5K6/vw2BTmKdBbDoM/tqsIYRZfXO3Fd/oQV1KDihY8P+GE04Ni1r5fKIwovb2loq
co9w26COwSK636OE3Dfm42bb3EWSHGn3nno71cTzUgcwnBSjzTCEQCh1SV0gIlPQNjepX26cQbDT
GAi8tN3HllWLdrurUqNn2y7IFhcRP7/OJapjBQ4RVP+tJ82pWCUJ3nq+AQyjLtsQc+W36B6Z4nCu
2FX4YDXRGPjLcojfHHSih7iiVXRNgWPNlivuV8XNpWiPaDneBv7uYmG2iO2k0GCRbLHCknoQJSeU
k0B7aAt5YKSjPpF6V1zwrRWkzxjyd7eyKvMiQr6yvaTVHcgaMGiHp1sXer5PAxEpA3Dv2vSrN45T
ZoErolZdYsMor9vrI5UFFO5Tga7qg6SjjZbxBNBo50lGavr3dZrSPxV/YHRDAQBqcgR+TKyM/1Cl
aDmESyHyzPFPrVHVfIwWaHWqBzlBLciQGFf4sZZRC1VH5DubjSQ98Ux0ByZh2gA8PtU/cXrIhHEf
r/8rQUVFZM5l6LvYL46Unhse7bmwcsQsX7HHI1dYaGuwT1nw3j2uSkk4JyehxK1llu0uOzWcL9fI
EFIB7h93URBp0Zt0MQ16z1Cw4pQm4qiDztY2B+yGXmzluVV6acPON0+xK4SYXJkV7/hgMQXMYLZA
WDuS9llqVYuCWoEQ0dH1GuyGqXu6EI6koQwcRXr9ub9yZVLLYyTMnTH9jFFgu8qSjLxmCJRpT2Jk
kzB2EQBtePFFGRIYOsrXJWJuNAEVOG+zzjl+/UCqYMtASV/kbSGMQzZ8Qcz0Igb9AfEcaOkcpYYQ
UfjHhY3QS5Be0MClTNGEbf+qe5w9kNwVy7Wpsi7gIzrpv/KQP4hXYcCI/bCo7WWR0onwWv/pMIw9
nn0152hOOEXgOQih85HKsR2sS/mQa+3kCoSTajci2ZjBgUMOhfJXInleowo3QpGtiep6GhxpxDkS
z+cRiVb4Gnfhcdk4jrHNiUMNzczDYiHr8gsbWIAoaX8Oz/zB8uGBSdY7/FYCg4lmh4bAogQ9c+mr
Z/ezuoZoGm2aqodWWVnCANc31u5Y1rbkcmAqbJ8bz1oyFEkkoRdDQMqyWCjsfv3gyuwU1BZM4Ofa
qbS1jp1t6MV6rsswo9KclP7VpEkRhzsDwYsQItcmcA14h22siw/+HA5Vlw7LT+Eqv/Rx6cfTovw8
h1K+SeznA+wXdLtkLtav7v8Ca7L4Vpxyp6cSPlOO3rbofSo/2+v2KcNMrGHVS9Qk0E6iSm1nqX9N
JhdHZJKQofERakqekRVly+yUAuvq+WLwNajv+2aSn7fQCFoqwPSc9gTG8/CKfxNUbL9mYngOIjSS
ScsjkE9EcI/TaOiqDWIt8Gxxj7LE6hbQ2q3vazhM2nad3XDK3svGLS54e3BnK10jYo0mZXb0CHBf
ASDSkeynv/o41zyQoezu0Zo6s6q+vKw9ZSymjP7gtHCxUXCCcEgGLA13ZaK2B3DoUocCG22Ksjy5
Ql6yuzre7sr15f/Ew7fEvAiyqhbXq+toIPahVWXcOW7TOJvMed6MZSTrywFo9+sdvhhn7KFWBRRh
/lIXiZzEBIJbXdBcj14PYfqenoLa5UDQraBX84B7obR4DynMpeTNJnDUGyrLnTG6JBrszGQxsdIQ
8aXATwhwivDrn/3OfgdUjolS9Hpv0HpPYYdoo8eWfcGPPAhUb0gf1M8OQg1GnCFNW2TSMsAE7xgW
y6su6r6WXRCTNYH3x+tGUP/gAAgO3v0moCePLc6xLU8Sr7KH82i5nAny0SR6F6dForXnJyw+5AOt
u3aRC0dMmV/84ywsOHfHm7aeIw+v1kouIakIWmwPZMyybjT3oIOTXeBMUgyEYQ4Ja62FZzVWBUkw
ta//25qU2WJKklv4NFQ9LEMGPUtwlZv0sa/OD1pIHVAjKi9wcS8Mb+AG7aN1NAAIKke8PF5CC9CI
AXDEp7stUToD4YXRwCE0G+u1LLus1PEgLQaGnSyCVCEHrADinfAb1fQoBGUiQVclouvWFtwy6BS7
MvRL7nbxdJZvTWzXpHrXhHRR5FiyDZmCYzDSvLcF/ckcyYu+b+yYoNY4QLu3hIM5s8Czqbps8Cgg
WerxpP91FLb2+920DNU9asKBfv5y7SXwI/gwet2aMhgid3YhekpG4PTiMzd3xo5icbX3ADrUmb9s
7zhN5Jxs8iS/6L3taFuPCy10cko3uwwe/s2AMVslrMB24vHUzXsaVz0tKflaSVjrcI8PQoQYJKDj
Cx0EwCy33WRpYkkPAX20pbHE3jLhb48NKed4DqGmirAHkxkZXgPap25LEEsAvUnRWmj5DOV/S8Uw
Ft/EZdiL/fcoV7Qv5uaqTiGMTwravJPfr5XIkLjBkH/NSRFh+jYqBAAE+JL0rZPmHSJpDcT858MV
onYfCuSiO3V1owc0zbrY8EjTuydAGg4NJJ4bzT1H/w3NjCN5Ufk2O6OpW+Z2pYi3HRJzZwJCLDKA
ef+vOmzqKU3wj4KIzS6fJvlaQh2kNK0LF8yMw3qg1uBqSswmzDOCwmT7VPkkUBprIppvlMy+4do5
x/ny2v2Ng28UP+awBhpPOi8l1RWLFdbQ6v6xfJiPNlp3bIpsP8Un8rqHXG+EaQJdHA5r+IM34VOJ
eLecwKE9pjuo6wW7uNHRDzkThtFePvL6ru8M+DeZSIEdk9InsVTABzTc9MgXWevbSplC5mcyh6KB
KC2rHU1ysDDxWyuNh7YlSUvwJIfqPWVRXp3nD12H9t12q1S12ZMRlqKTbhEbc+K8J/AWGb3rMDWx
qVoAqWhWZbMWnXJ5a/DAbu8YH3lcxBhuHcjraIZLCvqLe3J5t+ow2zCSv5DV72+Qomu8ICg28v+O
4LN3l/Ej9nw0PMQ83tf/bo8QS/ge53Sv/eAdd5KVlUp65BOnFntOmo4BzDu0bxa6DZs2SA10Yl/z
CtCGu/ZAKNJrMlkvwneWmwWtphTnRxGP/15FAUA7V/l+o8daaTXiCSlcWmdl35z2cMtbjWsTyN9X
MnA7TDdDjS8dwzFQivMjVxm1zRWVXvihzdIj2X7erNDiXkmJl9LwkbAoSF0kATFolJv42NNOJqpx
CHjTu/e2ERZmAZd4WrekBp3kIbR1TecPlKNbhzLXwWPXGWycLKFDpkBq13v9ViTYhRvaVetZsHZt
183wWfxccjerdH7BPvIEOdDBFWu4UxUsb/Q1LZuZvnf5y6SdzliiQtmxIx7YbJRb3kX0Pt2qSfFd
M94e/WP9mpT4/cCOYb+JSRaXEDkN8CjbTxHnohcjJCU1dw16nLdLX3j2nh/Dnt2YzUsmZWFM0nO3
f2Evre/mc0krs/+qqbCgZfVOujwEWeTPfPPi2l5nKKNNSIMbSDZ9oxvOoIs6PHP5I7uzW2ojXmmL
F9Z4d1x9nC3igCxgWO4dY49DZTxNZ0i4HfI2qgFR0H+nXRhL8X/nXlbDgWu3Gcmny64hBrYHgzwm
Joo0edCrMJuSKEf49yNshFbnarerCC45cPRNBOp7kontQ0I7pcmET43nXQduk+CznAbdxpo9VoAW
nJkYdJiVsurOATA2d+vMFpLctBaAR0Um8MX3NKb385zqXEOX4HFDKX7mjUNDhLpWEA9FDBQJgcuS
4mIK2JEpL05JeByq2OCFc8VbLfnNywewrCMH1d7a21vutUtf9UJRgmLxRpRlsR3cq/b23oxawk1q
zPE+7BL/4zPkbffiWzyjIP00BnMYCydECKHwzbpZoO7+jhX538IrOwNr2XifvN/l5xdgAyBD0VKp
YNhzlZBLvWeIBNTdhybv8f3GIws26rDAr3PBAQ7wdiWHHnmmYq9bj5wfF4/9Tx4hfxj07d07BArj
5JPuDWHaDOGb9E7VfIhnc4+RycV/3hMoqL2kLwa9isZe6NJ0kgx9mjX2Zc5/6AJss/yTcg8p9tVA
OB+n4DXxo7Fa9SLdVyZOcbAjf1q4zT1lToe92Kp19Ow/qL2UzgsLcy15eSjkhS40wvLKe6Vyc3eY
ugxN3d2lHLUEhSKhkDlB8QxpCUHzVIlhxXgCCnMfFZ3e4vAgbP50pNGd7ccOFSZDOd72gJxgnUPy
2cXB73Hg9dRV2gtN2jvFHZ0fij0MpXslObM9o4pSUIKWMADKOA/mZWm4YUNsChssLE4RT+6sHZNC
EYSKIozO4euDqRqDbGTeMrTYTAxXGHysuekSemztT34d7XrwKGvb/fE09MU/h0xu0w9CZ9uBXPZu
zDIpcZhhwSnaGQyyCKrqZqtvd4T+V3AvSHmbDSy34U+qdXOYxz29lEgAy+NoR7ec4zTIfgyLIr1q
br+axVAVAifr4CIoZZtadfCpXFb4IYqiXO44iYSPchI+SuSipfdeT4b6gurYoiq0Kh15o2AJHWP6
XTirhHxhpTWjtHI3dgM+IyVcw74pBVkaGVwXVEZ4ys/pbExg2c0OsoNsb6mbWtADZPQzbeH4RlwF
yl0/RfJ6YGxxH4uaAQEhR8qvxE5XrDCgrWlv0EqaTDc/slPFod5Bt5fLD/S/L/ZnGVJp4DN+Cdet
sONTwnCPx4gwzEHnnLkjtrEMpHgkOhdM9kiouMfdl/8eGzwMAQEc8lpfyHKwRdPfKz969lVAZoqr
ofWfTLXzQdzMzb3jz/9wieOGIvQys2Fu9N36eR2ytjX8NLWvOUYcnYxWxgha1pEl6cdh9iz/Z2pY
zlk4bIbYKBhqtCKGtGPvg0xUNyPmyDOgrtztZsAl021vuasezWgX9URfxi+OvLco+VHYesZOt08n
JC+A+JAdrn7HX1Sht2HaVwem6YtX5FOowjhPSb0nMzTnHOWW0W5y/+kklE+8ygmV4Ye1qT3VwF6g
muXboNORQTFeHuNQao2esjY7rqdUWN61jmyNGiEapVeLTmLhOnZZuc5JIxpnp+ftE1wgI84qaHv+
unQ1RfXptq9WUQM6jUcljCaWvdcW5oT2uMmjMwzFS/i9poFGvFQO+pY441dlf8xHA1SzRgQRsakC
6pWF52jVqtOr9WA4GxozFCFGlKDIX+L87Tt2j13216vEr2elFaiYUiMX3QnoHEN+vA4dgdd2Jzq+
w6QSLfTyiilCyaTjkrchdvDo3vByJxTZSiF9vy/TtAlqcDSrafkQyjpfP6r4HeaGdxUW7lK5kO4T
EJeRSL23P3Gpu0N+/ZOUrUDSJKoY5ALFTq5bxnntutLhtrClRZmtOQIFNvtWgRD3ASImR8UFAn1R
9Nt7tGfhA/T4suecQaLSAms65qBg5gQFoEkOVb1C8IdxyittM6B2XYryIVNyeR6MNCx0ojWRokHB
wt9t/5eMLkuAF9syXZKdgYOsNQ593ea0gBDs/qhEMV4lPz6ZLSzk4r9oLFEk5RyT014UWtLSgVae
YT4hrHDgEK0708u3k5wQ1JMn9X1GnYJyk5nuGxDUqUhlDAlVwDhhzTJjU9rpfXJU2guFdsqwwsoZ
b6NUwcU4gqi/nu0v2UUYHBvquXSw3iGSyYJPt6IS9iaMXCN2ABtfGN7mRKgoIa57SWpDXBRZObbg
si6hHFxleJ4KLNti0YEijtaZyaVc1yAEERqq17e8i8L+M4Yml58Dl3u9k+BLBdAscFcmm8c+E7KX
fpJ2i76RL57SLuGBIghHoICIxM8clsSIotEUbIupsloaGMJc/LXhbzvLaZR4V+pZReUKbN03PP4R
IY4OMs1UMeosH4MD5Kb+wzR8EY2fGDpT9qhBPe6rgeCnuYRdLjEO5YlAY4sEj3fpc9GwDDgroFu4
Rf8hd17Z46K+OpPP3XPX8KytZHHaYd/xCzsd6UwWbq49P55p0h1RVd6eXyqG9qOvyl4BqHI8Bfcx
vFvTqT8s4BOK26jvG2CLL7oKY/ebGfEg0ha1OCQXb3OTXuh1HYV2Xv+GhfiH5o8xS3PkyspNGc48
gloC9jtbmLW4XNtS389AIQH5NUam92ZTEnr36YMgauFcsWUc8X/PzZb/iDfQzVKGLae5gxFS2Ps0
ISGxCt9W3aP9TinKxDKwE0EjwKBKBpwMcLSYZSh53pFQ6M7XkiRrzkVRz3bJ+QjxkvqZ1TqgH8AA
VEiTCWjIHuniS7zuWXRuZIeknpr02XoNYvTIWXiVsVuGH5/qCTRjv8juE54arFETYH1A3bKXjigO
XvAqU+Uf6fIaw1mGIHICkNarkUGWBLpPTnFLDofR+eZM5L9R7D0s2JgodsEzsxUNXRpeykaU/WBi
oFEu02QRnIHqld6bU1D7/rUKTELQhoxpYZcGhwJVFN2p4ucS6JQrREw4fCryGXhOIgTAGw53zmXt
BaE85MuL7m41owqQAXFLm5Z118+GZVojBka0VDExxuYX2ruVUNTT2ShZd3C1pBZnBte2SeKXORfi
MgNduq6dNKyQ5Nk8ndsnzCjo14pbQ4UFlBn6yrIi3Bv4mY9qyY/jyk41eE0/BtzLdH3QXfTvlLz9
1oqD6MRoCeomBejQQy0ef+UcYcZUWpwN/oxUu4TkyYtHKCbyMAIBtsNEhoq6B7o7IWtZewPafRhR
4i2gRUxzC8us6LxTH/GCr0kUOz4SAKLkIazPDXDd1FZMkGaP+V6n9rNIJaBu/OTfIeICkAVsIU8l
WBAxmb0yidu5mpv+z4VVgHbSob1fe/x52HdFg9E9qtKhAiwr5bS0VSPNK3KMg97McofLIbCw7yDS
YE8ZtIQugfUL4DV2fBHazCb1UJsvT0vkZyw/TNMru8rapJE8rhk084HznjxC4Q5LpsQEha81nNM9
M0H7/TdwSGkhAIL9JgXZOvnWash7FYLMXmbYqapghOu2awV+2UdgbVWt5D41Qeyv40AGYwL5RrVF
aCIUpj+uZ/eQfRwAJ+atvG1WhYWqsHdHzyl/PqJdsdvizhTfrkVyHyS49KdF3sMMR76l6pJHUjy+
4u5FYULwTduWmR5ZV5QkCORN42msshD3+GU8UJu73Nmvsx3VwdWcaEv+7lC/l3CCvA1mX0d5KBLS
/osUfVigShSQea6neJNAPv2rT3UXNqmoKgR5W+Yq7JKOGgO5cKpjalMwvhdU48S5i4u1YMhfRQ/R
b2MEZbrZaErk5HcEZ7Y/w8yGi1qlaRDFugYIZNnF9OUabdePgODVlS5CG4ZWKdBU82Oqc2djYsQ5
0bfjiUrHOmBTIfGpw9rx+3I5zvB6z/XsyY2SZEvKYqGLsL9+C9DPgpgxw0JVA4QjRSIIDFjiShCg
jLoW3Dk4C92R6L1MKX4jSoOoNeDgpybJO/dKo8F37p07Y4aa9SN1ZsYiCGiDCNnUVSlQG5pBkdyw
mz/UlDXTbzeSpjT0eCBY2R+5l0SLd2XjLrBKsRgMeXrULuza6AjC6x4gjGp2Qp2StmevQJfeFAMU
I1Haiq6RAZ30AkifaU1hZnfLQAcewck9B7oTs/NMTBAkC/xHuNuz7Pysp48TzjVuK1rbCVsHt9cv
NVX+suuhKKe2VfR+a0MHkqSBU1xDifHRKNVgE1ZvYI+ZlL6VAXxnJX5hSzlz/27FNSE3vdPTyoQX
G+uIluWL+8rki8QH5hsN8vEmWFLFGN7q5ts5ypxU1dJwA0pTMWOlFAMTg2E7qtuhbszCyWsRmXnf
7FYb1XToY0x5hB+njrZSpsHYSK4vMQfaU3W9VYafx3GBgooIZF/i461leWXak9Ydwm2NYMKSUKeH
0NuyY58/C2mPyF+5cqzIjKe1uBKaKz3SrE3+7uT3r3eCUWXJSTGBkn0V5tFYYDMAgmqWwLL3j4uB
BKz+X4c6CCopRCpPOZuQmRqM4qlJco6i2e+h/Ad1RDijKoFaiEfNTz90u5HDPYuUPIrC247+50Ni
Qt4UwbJSNXH8skekf3LrBSvg4TlakiMH9S1+U7igmLBt7rrMKG3iKEiiNXElG4ubeTpJT4UrqbB/
7c08+lZkDBR/ok57OOS0qDgo5yHySiVsaFtKeXREmJgUfqhKiuHcOkwO1yr5Y9yI0coIiSXhYOgh
qAu/BHwYpLj0E3F8OOA8oZkmjExSPeimQr/i2DIov0blmxXZveyF1IZqzW8frAdXWBqVcJhhSfm+
0YzOhlU6/E2eAIACtGZ3oN1I4GlT3AaQXNbiUsbdhFldaNPkSbChlvvc+MwV4wGNJ5tLWDf1vM2c
BWcwOBXYdlN1FYFQEDRK+OeUfnZmHAdypwAnlqtskWrvE5oNmWGSHoUHBq9psys72WmJZAZGs1wK
+mncIVGHFE5BXK5gSY+R0jNNae8xrfammg/3g4iBJP8Q1NMcNF7hdL56OQ9oXVxaA9ATCWBFHMhN
nSH3hJvN9O/MLEATIPF0ON4SVHUVdYGLnvXiXacauRF8Iv/XIBzbZb/NjzmrjNtcENlqugN4XKYW
wSj8R3kDiXolypPx2slMpaK2Nbt1x7P0A+oNHiJLpFdhkkNERNzFm+jATw4ZmR3CCUQWL9jRudQJ
lkb5n9ayNXy3FI1LbAkQr4bJ3xHVtLnP3iCwZRUpL2mWv67nrykHQYOq2R5E5S1GiPQ0AQ0YaH7X
jF95lo/uwqK/49PMDFcUJm9fgHXXvTfPIuZS4GhML4DTX2CU8EOBjzchDNXR7DR+/HdWCpSFQd3z
hCdLvqNZJU0pFOvxYB+Qv8J6bTot2Ga/wTKzMKx2MEFG7esBuzURDyQeQlWrh+NVkgWxAK5K7Bty
TCPiijY+dYM7K8tfvs9oNeKd0xpTlTUlPBxrQF9FQDB58H3R8Xk0C6/soiGzJDEHaN1avl6YFMyz
KF7j8D3G6IWMwh/ENXHfi7REPhGZIhEMV1T/qi3UMpPbKvdQamHV73nTk+GM06E9neucJJRdS72f
ywyyv8JQr/yJhWRtUUGCeKw56GyPoBV33DHrLqIx0EpcDnjy4rZ43ztwJNReFgfU/7WEcdg9iFIv
TsUBpUpNZYZdORTkaORq8Q7YzqMFC7MX/lbcOyZaIDNZxtcSAYWNcC6lj6qWFZZg12IQDcTV2mVK
7mFgnSozh6LhynBUxdEll2LxwhDJChMzok2+7dRMS8slWs88geFXN2k1bLArDPagOS2hMyPPrbop
cNDETPdsu0+2czTAMhQf+SvSfYHG2i9whZORLDlJFsnEkMShATdD+xGOXKZQ/iMYArMrmnlEVAum
3cwAMFWEVFcvPyJgQKyg589RYrHcKr5ffhzThvQ7v+3dlu3fKOAVP0uq33WgI0o3syb32HIPMoQ+
jnzeBOwVUpWFqYv0vGSNrtajIgZpB49IHuzHUoAQhVPUh9ln/BwiX3swZvFL3PDKQSYgODOj3woM
zwiOLB9ec972C2Oto0lUrQ7ICYiQws6BzgCOQGhs99nnfCg66pQbi9/i8Awy2MZ+eQyXr7OTzKi+
re2rcols11ozM8pvcvGeP9H+VaDYGhiFzj540SO/tngwNvEvCfcTql2pbzRW1FvMLB/+aMYMjcMO
1x0YpAa8g7Jcdtn7ou5v27GmCVm4H3ZHmEe8LHRkXPdMIws52LaG7p5cTipkKPgTDTr9xqZmkHCJ
kT69gKHI6Z8NH521G35kHwjVhxpMnNDheKQEG7VgZqvRYfRXy+jUh6lO+mYt1w9WVM58A1yUhRnB
1LfVYkERIFJx+AcNprAl9Cn09+lC3236H0ZzGCrq7bBNG0lthXP6MVdBqdloaVOx9tFFR5pGPcGe
Df/aHq/rKMhsQ7B5AioS69Wz0HFzY2YShpmTYN8xIZosm/eCN0LyVNybSiuEWGdSr20HwPaCvvit
xZQilnW2aLHKBLFMq46mxkyMNlFGE7Cxw+RpF8pa/7VCtEgcQajQSKGLkHYqoJFlCMdzYwCus6oe
b8eeQy/Jc6qtMyEsDfv2jIJhsd+kACrLwmmyDmdHUC95Zdbdv84WRg1N/buH0eN8DPL6bJcb0Yxy
8X5bCOXfAXPVCfcchO8BvHWmMpgfCXjJ5mp0QRs5r8PhYXTVFicAy9lk6FZxzi7yYkgtK1+6q5gK
tyKqGym3bDt99qprPiBQ9poTyE+i9AZQD/S7jNmMffzmzaMkMqyG5blYT3j8cOzXcbV+oFjwiMVe
WrSLzEPwAVAmgVckIGVXTM4ve3HfJC5FN6KgGVmDLWdlSMbJyY/8YQNx/SBPONrwN5Jnh3lhi81b
HnXpIsNYq7R5rFwTcOBavwbenBZ/jRIdfifblbq641XATcErFu4uhyi697qKGySe6n8J0OVbGzZU
mOXjvo85S42kw3V3AJeQKuqEpvHTd8c1fFbNDjeHzy9giQNyfx78rrpf2HawZqq9Nn33p2NW5q3m
BmRrYqi26gg57pOGFOIR+/Vi8nSPqubPJuC5vwJ9M1oXEWQywQ7YxaMdaG0c8js4J8omSYXmHelB
kLLZNwNxgbYs9d2nTPr7z3Q9XEVP9iAU/hagtFbtiZX4biBYht+vIz1/+55aSVOem4vandSnv6rr
zw6nyhoDXNC5RIg6LpddzEdeav4sLnMv1kR0d8Us856STpThxwAWGLMwE9Y5a5LKyQzxdarvjYZa
poCPAWLbLNxFry3JDub+Xv36mRnqgcPfULHVB4QBv4OLM9At3fPbScpvHCIGURPuowK7umb1Tki4
R5CslLIwRF5R/yrKDnL99FyxB7s9dqxZXrNhlhqF6ADXnI/FegHMCCJ5xNiafF/Gbfggqm4wF6KI
cjWnF9B1NQBe+8HVpqThnJ/ux1F2+3uC8HnoPa5QmTox+y35r9smj7roYWhdapUne/Wytv2KOwaG
gt2nYsTJ/EpGDbBjroky5n3DSCEyZV2ZL7pE959qZz7RUBPAevjxINFe58w4OJ+GMYP6/7hUQgXQ
S7rfIWG7+ZclcDvfor3IqUrqVAj/IUx5nZDAb8zQCdFjEqK0v/hQVkBluehPCgJiPR3SR2Op9w4U
i0ozbCnFedl00fFyrPB8y1ILBxRxIDe3VRedIQspmiQRAjzk1V/UezQXhR+dmsrwLMifHVp664PF
n0lWoHPHWFYN9DCLL/i6KEXG+RG1aafIS715O6gXEofhhI0FYeq0sEYNt560UihzX1cYEO92xIdR
MkIV32CfYTfIfV8svXipj57eKYpADHulBqHhZvW2kBocdPG8cl36coebBCmVWQ9+dydi6PGv3kON
71F5wTZ/W+uav5KCQJA+JXOe0Cwcoz6jZuCaXtIM5vbYh/CYsQIo6AN/PSW7NYOIJL5KKAIbgHVL
Br+oKnqj9/fZqCMM6CirVB6QZCYjz01FV5gsSYXC6gAt1JbD3CpEsuKBpDx6OJVyJKGgJkk0BtpA
1p4ydBxg5ZxbbBtiaCRHT4CWrDzzalaLWdXpdQpdX6rGr8EjsRwGrJpk3lsu2JNFE6PjEYvartJ7
bQhQJKJ1wn/UOXwVvhltCwUYfU6Bc2I5bui0Ek+rzRqK2ffQeXGtdwEmuhZidnrBpizDxpfKLAP6
LpkRzSt1UfDVGHIQFYDouqm83ae3jl8VjKOBeoDLWy6RICgCAuPduT31VGW1/7OSFFMrS4TWYWJL
NxStn+tsOZCoib9sW0lGC3MNYONZ5VDuEIvJhhklG2Ejmwdxl96PSNLNnb+XoozUdfAWyhdLyg3d
C1N0AAEOmUSYH3UIW1pFnYg+MdIFVZymmbEHEeYtZtdK5B13DKUVEkYNoPWDqKvfBlJPLQESp8b5
3IJQULymT74LZCd9wzEsBBgeAnru6tc/VDfKhVtraE+h3KxB00Trvan3TSvHQafAsKtx5T3vjVAS
tTRpOaoSpEcIO0evvxJuYJsqnSWxz1WDtaZSmax7MeHO5hR6TkjV6Nd1ncVyahVePyp4AQ/xGnlJ
2QUe8ovTv0572Z1WVm9zRjZWATRrMrJxeZGzlbOJ2aFkFvO1tYY01nqz6Us0ujAAWNJJ6qTywXdH
4P7UfR+EtgkK0zjMzHKFyVCc4P+vxV8sXgPegz73qTPPeTWXOTSclUVwOGOtLmoMYtGUWkYmYUF8
gSs5h5J1EpggFCvg07hMhpYEE/xZsD+Wwq7Z1acoYNr1FfqCB09V8u3WOuXwMGBq1miAGQAHK01s
k47E7evUkvCGteNV4PzZIUKxmCwVl2iRfpRR2n0ke+LnrDRMIx05KZHU2CFriaLx13N4Ggud0YhK
cYgN2B82ISV4HCR3k+hEx2Xecq5adQ9HsYkSILCCd31QgFE1aqP1Kbb0Wn/70sVlkbOIghFus77i
OIyl4sjShajyBOyANVhF8dsdY+HNFTNxGpI4PvLWdg20ykoryjXg6BQqdWmvXAyjLKEB3r9Rs9Mg
uwr/t+EDGLp2cOX038hFFIpK3bfurvTRruko/O1LnD0uudbH+xxQiy3+UzaN7BfIcNYshp4IzNcM
E4j9HkPDiyvIoGQdx/DUhDx3MpmBTjS6RIYZHQLASAzHormkKC4G+p4+k0anLZ1kPFmvuyCYAzVa
WETVXFNvjoN4fcAudIZHOp9fik+Wwvmawh22wsxHTHdJzxQWVyn+GewXMAooudRyUFClocdOB9wG
XbBh8cLWlyDNRjU2k/exzkEfg6Oaxe82f/8id0nSS3csgre7wAcxhPsdoCQNvwq9LJD/h8O8dsTy
wth09LtjjB5w2wGlXxTKlCIgK+oUC+Nvc9G4rBlFIKSKPUOuckfTMmKt4JvAm4IYZv5dHI2EMfLp
DqEVesH21yuwin0lZjbEtsDH/TdAdGoxpn8ScDC9q7vTGkcrnVPxIrCZo3NRZ0ThCjPqAGULOBUh
j97H7UiGzbfq7QuR5uCutXflPdmPn0qXla4LAy5HeGE6aGJ/nlyPMexQz04K0Bd1PyiqK7L04Zn/
cwfzDyFplcvvPbtVds6ZbU2xVlUV/JSuMoBfili/dEJP+xKaE9ZC9EU3X2veMcBIzGqbhpakpxVu
3D84wV6EicjVD3IeWydzgQQZ/b1EPiZCYr93nMIKYYiL9GSDkJS3e8Odrj83eFLOXUzmZuI4w/vL
jcdPu+Duj+qgWiTEpawLaMlisc4nY0y75XOs8pl2jh9wqEBTrkS52xAbpFiXsca1AOuKeBo/2SDF
V94h0zeW+yo+VKalygLx6H6kUAFXuFDBurl1wbxEZBUHAg3A/jPIFPATxCXOKwSru3B279aSt4EJ
GrP7HZvOq3khNbrX5g3AxYaEwfYqfKt0iKbldx5vVXhdnDb64rXnpb5wv3qBYdT5bZ+DZHDgn9lI
pWCT4OJlhXu3R/dvm+NqSrpdfGSeqdW1FCaSBzHkKXU6D5EusgX05v883/dws/R+XuTT8IFohZCr
c1p1AEc24BiVvmLhLFaFSIkA7pbY4UIDlSYRlC1NYHO2xdWiGjocOlf4wflYgyZTA+L0010iL55g
J253bSlM42LJBxucqT2C5oUuB2/gmaAURyy0Tt/cQrulamcbECbbAahf6RhAhrDo6DjLSdL62XFl
VYNjNZD07g2rC08Ui6dsNIDud4vE3WknM9+SqbhNeLGbrGikWTD38r3zCFox6PojclZJdIu1ujj8
Vlpp920TOfrPc5wJpvFJ3TUYGRr4phdSgF8FxfuFKZavXi9mF7DvNkCLDVjt7g6J2HqFKQPYCFrI
N3m349Cd+xTLbKgS5ao3zZbqg7/97Ow4bxNyPv6joiykLiBcJIErUXFcO0c/t+4Tu67a9S+zvadx
XqCvr2pz9lPbHRx0oF6UfwE6e+26deM7I9hcYQzO2PiO/Y2mjYKHG65agjnSRV81Rs2QYaDrVo+O
WshEZ+8DeKHy2RNqtbhnWt8HG/XjNTmd3hL+Lqgn6o7IKXi9Ud7hSyXh3ML3jpmU/hxt6ACKNofu
fpdTxtHQTrJBwSGNtNekJhLTP8s2hDMCR3atbhRMnqBcEdAE4UJa62CBagP3SkgqkuO7ngBTbp9O
QMc/60ZZ0QvAHV9ijArEsnPhlzqAvQ8jqsI1zNIpQ8W/I3A8BcUvDxKm4clpWai97jl241NEzOoP
7qptw2LDZKlkw+sveCT4gQcl8gakUIYX26OZRCrvKqfoWhjZmIWQuGeaRHt/1gQ6t59cOw3SPqT6
RIZLcGsJj5bDnzjW6ug/JjoC8d+AGG84ZC3VR1NTKku1xyhf8d8K/mmBlluAl+Encmu043epxusC
uclHT61o1ZPSAmaVIR3RrVa80Yzkq8/hKCqOT+RLtBt9plemz1xwFsfZVKZxV1VsI/CrzZDi2h0u
l7ox2NBhD+0J94Hw4STbl8F9GIwqaQ31pkzKKIl8KjFhcs+wt00XAPg38lwpjWxzN5OdSoJNgdA9
7zQSRV439ZCeZaa3fH6WmsEemU4jouBWr9ygV3h9zr4zxgsQo4uhH6FGXAwTZn2fG/lAo8Pe6ppA
IhLWOcmyJIls7uZSdOMjwiT/VW64UBI8Sx3K60fAksNIhenp9pAsoqj5Y/I4BeA6230kzFXMEyrn
d39zl4KtcuiBZZ+OKh1RHFFRx5xOmCVQPeH30RUdhhWUvu7wYI0D2KpbqBwOy1cBF/PjPd6pH1Y/
WhgHMXkdUadcP6cuw6l4C5O0c+IoM3ADHpywgTDi3HPqSnbidnz+BQJ68MVDFG7Vg8AEfe56EijE
cNnuBw3VAzJfy6SsM0mVFsr0a0+DqwbnppHSU/ean94FCAXPWde9PLKqddYCS6TBq/j2ooY0IMUX
oz2iJTvPF2OzFjmSGr/vt8/y5dj4f0fMW7UneOPN9NKTgMkzwIG3HK6G+24Unvh/MVp+KSxg29YE
hiZZGTj1PzHF6K+/NE8YFvBJcLY2iQzN4saOGkdIM9P6t5IpLXMCGbwlnEFTtURp2gLdqzryx3zE
ky66vUlM4bYAFHh8/RMVtVgxuuRoQzanEwoM3B9qQHIFJc+2hXcL8FmFDP8SdFEGjkv0v/c2apSM
QVxoI2hdzQPmd3dS37MRMwJsgX8z31Ybpaaxh8m7BsrPbAerzCFXBh6AHYgyfjejIRJFHmGaWNj3
ximMdjNx7qvJuwSVKj2oH0wgosgPYLuK7SdHab2oX/0KTu97cgUGfcEOQoDjHhnJZQglQtV9Se4+
7LCShnakazNwk6xOn7Fb7a4XmEviHSWwgtfaCrVHsjFfwt6kYlNYc9J0FJvYiHliW9neBR/iGoEQ
ed6g8IAQqsvw3o2ml7R+BQVO8CNTbr5Y+KYgB/2iPdtCc7OchDoZSfEm1f5FA2jtibBoTiVAdnZ0
Yp0f1YoYyUjxExsh/WR/rbKwHlwCsuY+JRwVaSv89St2OhBwF1UxLsI6bvoatwCM/PtWkyhDH5wB
t0CsSoQw87MXG0hy0yEbOADHjNsIFKyyUCmZd4aCR/kXZMaLbDnMgDddhrBEfmfzuZLb+PSGbTrl
ANqe+3QiP8GY2t0UQwIuTFcCR+7Ce7yAJruOqIwQJ/OLQwJ4Ry2kUM8+hI8QrAEzbxL+Sz9PSwlS
18sXEBfqd97kS0RjqnOoTKX3VB2eLBYbq8mN7Te6HEWn/rdDXMUPnqHmAuR0WNhBQRGU8cSQSNoG
3tzedrajAvpCT/sDg/zn3b2mSSoOk/au+9FLpl24ptecSg4A0m/FJ3vcmObm8n342/dPXt6XYmqN
QXfb/BE4wUVo8SKpLy6qaKyjbT3eYpfFw7NMxlg1/nLFu/4y15izBiSNWYDAGmcIDVh1fhD1W+lR
WyPApQsf9neR1lnB+gJQjojO40MX2dRr6+/jd/9EhtqGQJ0XlPWSTETbYybi/VloB9m4pbJ+/R8Y
xR8P3L17vgwP0gMOF4XoLQwfiYy20uktHOLanxWRLDiQg2T2/rmUBUuROCzMxlQSyeC2ylzag1r6
Rl/73aqG7ieQqVYn0X/+b1nb09/UTfLJUJTdxWffQJIKVJJAUo+fjILvVUourThreaR7atbiPb6x
sPkApq6rOFMKzDvtADIjQlC+kpxAxfPloTLeP//s6UxAJ/R4YdZ+yprz7qhpdVcfsH12nANK3Pd8
+W6cdTvdI09LXA98YN0CLgRxmq7LkBoGc1wQfqdQDb2WZSA9xSkZIk5SC9yTZ9yPgv/6VY73hr0o
RWEEzG/cO0b4RAqEhPeA9ccqy7cMB3CIiaoEBtlxVNeaoN0JPShaFrb0lrkwW63FBiWz3j+hE4Vw
7DSXuzB+9NdUiqTkLGGWOivDuLljrrucpSbJ/EMoSa8sglz8vloF3hHXz9zQWaUYoI5rTkaE+uQM
t2n730bat/lqvzE68urTNiAZZNo9CxUix4jMBoEhD+eOk4NUh46ZwTPMW9wiWpPg5xHH/MdlzB57
IcN47LGvOyJgopz/2H+fTa0k/y4ItQp4RmYd1ql3ulaIrkOcAa+zzx9YKKWRLkO8Y+2NR5q/94TV
5QHQlIH5M9mb7+qwtuZga2XMZ5poB3KHDxOzWTzkgDNfqj5mqE5IHGo7vtUjXZhcid8527wsICDx
jnp58VHDefJWG5GTQr83h4dUNZuc88rWmY5yc+pbqbCyRcRCQkXAzRvvxjZOtIaYwXQpeBybu22R
KfybyUTFbWD1NVulygasSE95rdbY+XfwrhRFV4yIRMtzEIs8Zh8xDPY/1rsmShNVn6hIiMA7fRCx
gud+eTqIUQy1Lz/WZ+LdaVPBRRXEawN3G5NBzL4KY8em+0Il4OSEeOGk1BcZ8hFjR6UZopWYtb+k
vf4NjETbacI6ef+wzpvVyrlSjHl6MtzuwWwAidDf1llC5ev+VRq65Z7sYcQBOK2tV6MlriTA0dpV
kNI0HZJg5pW1YOyQMI4zXIbW7G3TfC9nFcCGJe3CGiN+6Nrwszw22lEg3LLxzlhRP5KFQZFbPqam
qkpOVGbwT+ZVQjCtC95FnCO8GkwLGHDh53nvg/xIYYsPnC/HOCcSyaSg1lEeB5fdSy54owmH0aw6
R5Uo2E2icC8uWANTCxn4yPxSF2LnYBjYzZPwlCbRSxyLFzEmjFMAbOr/HumKp4FM0uXR/IYnGlCY
ibPGHPOo+RkRft520tIoSFb8nNzqzCIyFjxvjkXyVdX9AocATN8jR6Mh2nYMyBAEegptiXuh5mFY
6boye/FJbJYyKFWpvwUJ6qwCXSZL0n5glteZN/O106kdz9U6Cvy3m5rv9zUWRCN/+Fm2HwK7jf7d
GWLWcaIpaDoUc4C/Kn6U0FY0Qb2fKlFt6WPRXp1GnJPMgMgTM3H7slL0JtWudlzLaTfABsPBWsH7
FZC2aZ39yC0U1ClMMNnFkVbwEtk1RKa24cX5e7Q44mWCDa9DXMQLoiQMj6flG/z9e//cHmJ4IEhW
6dJRef4kUko6JCBoobMELFFYVoYk/9pmF806LENyzBOl/2cauWWECvmPF5K6Ks5xBz/TpBeBe7pj
AFptgpgKdKoW3juY7TUEe/wVgbGd625a/UV9j9eaWb3s0+FamAqg0uq2hRxNPUkATY9UTBJqG3Bc
NAP6qnRh5WyGnZ4NOUan6J+bcdvv29jObzh7rw4edy+U6kujmHzeSq3Q0RLTbMF6+WBLaBYJdF+b
HIw8EVoFa4jdIiqHV/Bpl12RExR+RCGdXK4TAForkc0fK/yjGt+/ULBcgBTPTH+NbCBOj1NNuMP5
7ZATi2VCXqr5ig/WC3UckMz6xHGztZLmNOQYljNOoah9l00feh3E7Bm+DOS8K6ibVB3BvaqyKTDH
ScvdOREUt/ewLFJcCZ6L6PAuFrP6Eu44uoAlyRWb+HgLvsecWnLTHLJa8Xsqz4f9iJ9D/FIqqIXq
iMw2exs/MMJTl9JzjiJyoLi1zElpXEHeVtyhqsmVJx+nCBqm4qTchDy8AqFou2U+uP+kYDAlagNe
tCTdPMJUzIwRo1M95buhdYZ94EJWxNTtxbo3xOrtAB43zEq3DlvqOBzONu2aTPjRyHHuSXGx2AaG
VfrbYhDRUymKAl0oU8Cvs5WdwKLkTFSnkVZWp0XS67A5yykd8ISdOYLCihquTUAsvtf3DtJH63n0
/SjPguG9pr8AsxPR9zfktOOb/b1QE9sSHimXGl9cCdOouXOETVkhESTcIZllRYto80WLiHc0v//k
Vnu3eL+gBNi7MSN7psrfilYsepQOGMnBylLJX0wfPDIl0tb3p2ZG6xTszGgbwtR5fiN9KPqDe0V2
7Xz7kqgy1iVWjQdarbYr0AXv3bAD6Oi0ZdWUmIWLcY06yI870ii25M1GCrcZ4bBnnDRNB9fblont
s4Z4goYMdTC5utsu1z79CE/YDiBkqk5WpqvQYiljNX8tAr20lkAdAjDJMo7j1CjGV5v+Jcnojlpu
jDcUwS7+aOpnQLpeEBThRPMEHhe9e1fQDm4JKDtuwrHU4Oqs4pyoD66zlfh5+lukf3pgOFTxS1do
bnfNxdkG5N+XkVoBqRkecyr32bhQljd5ib+quQERqK1iysJSEhQ8x02ZbmHe/pg+e2KuZp2W9syH
Y6+iwuqaPLhK0KfBBVnA7ybEOLJDgShhFt9Qmho2FpZH7RpJtBB3zDOmTFbU+R59bs5VfDPi5/Z0
kZpdBVYELXm2cFEMn8SxAMXUHtcSGYWLtds+V2urtwfJdsZsEw9XGb9CQNlpmEBeE7ePG3KHkNPw
8f7M4CPEqoMAeV29B4JLaZnLi/L+44/QeKWwPAkwio6+p61uVIGlyJ7myAmCmZM5cf1to62QLNpu
PUDgpgNBgyNqERWrx8NfpDpB66JSV/hNZN8wY2Pj7cB24J/STLYrcYGUCioHd5xifV2ICtDzlLmN
r/0kZ4YawtwE5mdngssprwMVueFzsFWYnY/6gMJ6tPaRFK5KPM1ROp8Sj+j76PWNP+1c3Xwm0WTh
mx7Mt77EDCmZGQPAVYalgUplyluQqsIbIo8CDIWLYp3XpZU+7t5RudRS8/s+ZAfczqt/fYRYjR59
CSSTkSt5fxBCIxfp7t1oxSgIepF41vpNvBjYqmQ4JLWVMaS0+i2HQwmL5C1S9gPRIskhl/OBHHdZ
9YxvqspZfIceUazw1HtyvJYsmI1o2OBtWjKtM//g6xIa6WSki0ArFTyqVdX4yRu8m8hFENsd7Ehu
eVgopUHOfvEj9h//SkOCm79vgI2i+BNRpKX0CWM52+tSVIWY1AEMX8YnI8BfYyoqFOSlwwdLeqP5
Iytrz/Q/sbmFeKhjyTE6AoRM7UbONeULSX29U0ejHteV4YFc1x8wLUnLG1kdjP0r7p2N8uwcpkHr
IhF24cZmBWeNoJNkmy5Gu58hakqDJqiYfcbusV53MZ4R4kQsLC/88Xx81h6hoKnvqqQmvainUkR3
mzt+ktheV7sPFpZeGg6dLq8BH4CU+xkHUsyJUkGwewLmMIUYoDTyg19gZy1pn1OP9cDLWMX3hY82
9x5aCyW/viOcjkHPQG4SjG7YT+Lsi9dnLBXv/n6q7V9Me9URzbkLJGjv7087YKGzJjSNm9QabGDt
y69rj8YM+gTyrDQq/6sjOu4hCHns2D5zt2+K0ZG5MTT+HX12Wuj8RbLxAyAQIdWBt/n55I+kmQlq
fLZ/irDt6r7eI0tyS74dtVdvdedkHoVbTZYZUHAOiy7ijOMLnBhTkRH2jl/hw0C/hT4b9fiKeq1A
P2nxnDXxo+NFY8IUF0vpKtwx+jFLO4uYBNkmBVZsR354MjOtJQFsKaFfIfYtcn0qTySEN4mAaK1z
FPmCKvTUF0vI60/U6KPJceUnj/DVellISBxqmgZhx0FIvlZjpE15H3ZtSM9wQvAUKLix20arFBmR
yNhgMYNT1fnadEG4YofLleUzA6sDUL+dbGhteywB3s/P8UM6HtNmkSatEmaJ0DTEkaX9vkWuRlGc
v2ykuaJGYnQwtwALHHEh+z4kHG4gWPOCOv96zLTTBES6ss5LI6giZbL1xREq9e/2/odnBKlsuwgQ
ghMqw1fR2RjGbuCBIeknw+Z3giRjLYioirMw00aS50rxaQls2NwvaKH+HKombVg+bbdcfPrYCzNy
RBI/iHGNOuVJommwazcY8/OyAp2zaN4xcZeEntuspRLybmbvhze8e1k+10GrSTa7syWvsmwfBL5h
x2KVOqYDKYd3EiLfNhx+IaQ3XOAy3uEI2iClmIRVdXUlMQN8rbnHsIWnYX2ipv1rMvMl58lx5GJo
OlaS10ErAlby4CnrUGrR4z+adEuz306luKdxQy9Uztj23rDWhZv7RNd06QgwsEM73x9lJonSDf39
GZ3uCnNGDUyNGGYvRNOLOCABBdHeT5zDawxP6C7IJOAi5TlZISTepqSx1aZnqKVdQpETfmGD7B/8
51Arq+aZjSjKBKNzujjU9AFzrxwEmBD8GZ2oFIfcBwsUAlzJzskIP4ZYPMG7yXSWu6bIuCwGE0dg
pvuEAmLDYIK9BRE18m4095PhhI4gaIk05CcRhcktpf2pMlCsVWsr6Vg2CmZzKEISH7jeK2pFkK5I
GX1r7UEbPS6RPbO1G1+Ezc8j6cBX5FGQOEn4GiDHLeiv0qs/g6lIgg4dY2I9VH7vOHhDBEQfzvdH
UvshKa+AXitPNfxzJTrEJNzdddlmwyl9gWN53P6Fl7X6jDo9yTZE9tkXhyXuyxpWg4lJkfZYPwuR
TuJmDJAtSmwq+tlQGWWTWiIApv0lpa1nkQqJi1dalz1/vM5wub+0dupmCSdj/obrzt7rljLdlBUN
sRQAvb0CNzhvj2kyy2A2NVSeAWfDeIDfTC3ZyqezxSQS1485WVaNeSAiE0eZ3/dg3Tx7FkEl7X9C
aZDnc41lWfDVyhI+OGZLwaQVouDGm8NThz456YQKsIpR+UvTqsoYK7VE1url6txCC6HDkkvp7EEU
YyJc7O8A2cd73C78AzIzkRX33bvDl1tjjQ/94DHM8rUofmtNVfTJZBKifMbsrXos9Z/+YeX/8sOv
5W5PV9F73gyJG3miXi/l7W1DpFI4yeRDNeYhfjPwEPqDwxQ2Pp/5yvGr4Joy3vjhKDRTN8BFGnyy
1qcg+CAvhBXk+Cz5OWto1z/cglmPrnM9cnskbwgIGbf4aHLNarzZMtxmVDXC2UeCE7ObPTQaz6QK
gk9n3ySQwGMR7gLOaJ0NvPtGRVVNrWmMYUUY4mjP3zqfyv+4h8DB9tlPxrtGtMsyv+1VMfQbQeVJ
geHLhBIs194xetQMNXSwhVnl/gHFig8WhnmKBmupeOzrY2M7TqqxXWypKicG6mHj5FWdFF6LrvnT
EYWKoJSiqr4eUYcaPRcd+cLsLkCPpjS6OFDo25HMf8tcBByNcJF5iQbNSq/Z/TYr8GjaBKP+rTFD
oqilnIljeK1A9Ma+3GlguaLu8Ko2pnJPS2xV6OCwsOwVaCI+86sm1M4yIP3iYfN7baKlAimiP3eU
+wSRO26harmN0iZBSYpHWthmYwwO7mqrL4RAtlR5Wj52//uXL25Oj0lspDe0Ry/IBU3uI8P1GAA/
wPatFYX/TPDispBaa5qGX1Xg5AOt37mXo1EEbPIlpfFPOkbNVKJWQpJgJDNV8WFb/52eqnT8xLdB
5z/dvmTAcNNFSrdm+KV8xTVACv9TbB/KspgEc53/2Z8xmYX9vRsJtku15O1Uka5eANaauB5TnvVi
9hO7m4NsrJbp2CDkaBMaDcHX4XqGPMLjWdMYZpcwd5R1xV8kXgHgj7tF+FCEncYdlRJPENFGVQJP
NU88YmoE6FY+odA8y5ZI6d/HAWpcs7q0m4ElptlstlolLDaur51CzEkAUgsRRIqPbvlnlSGPPON6
5y3W4BkZZ+1kPaPdoa7KYRKdCZMO2u9E3vq7joXWUxN3DZOX3mmtdG6vgp9T4gS1UPwoupqYlABr
ojYfwBU1JwrBcuRHpAn3uyhPIhmiQBTaYYCPPaJLscMMaYEIlAOcQSsiZ616oc8E8XiXdBqg2zYN
BT708Ifd6YD0s9GHPxEyGcYAQj3/uHJoucqK8j8W9x8rLDizOp563KOkM/C9dC7mINDifvnsb4OE
VCjLbkj5AlhKQ7HTv3XrrEo/lzk0oZdy1lgpct4Qmflbg4hpkMxEQp5LNfZJ791QNRqERdx6UKk4
8EtSE6gmBg0bWpScrNKs3ctqTwLB+PasiqA6EhudC2CSdXO+zxtzlcza+V4KFW3VeDXokDEwFpNo
AdyHA2eLeHVPkxA+difyEE78rmyS2a2H0BojlHGYmas4bfHnDDkyhxQNxhHFMFZwjhHnoRcfFDPB
sogK9FDXdlRDX5VVthluuh+8Rl7hkrQCoRSpNWzehfifyOIb2LVialNPSmb6T3y5Bo01lf32yBM6
slFKSyDykFcLxIcJoT2/hfOROjx0YFs5QUudZeqf9+6J+s8WonP+VPpTUr6+XuT93Pm5s7tXh+qA
a5LVKrsRnqYi66NxRlj+/8OHamzxKiO4zH38SJVvAlM8Or69YNYoWR82UjeHVF8+CpGKmWdtVc28
rBG1VMbsfN5MAuhCpHI3UQqTuGkL/4ge92/9elnCsgNhuZ/YovtUXKsNHHwy8TIAIK0JNZoI+KZT
d9O1eKe2MAK4GB8bKslaaXtmWx99glAg4twO9qLME+Mw9l6ZNnsl0pBzcHDI/Px8E6mw/YWqaEKA
3ra3GUTrTW4Kdrunak2huk/8Y0vAD/+1DWtYkoAFjqQjp1IHHQfsSvWJUZdoDMT9ACnZlD7hEC6p
Y2CX/5KtBVqPH847ndLN3/7G8Um5BYUj5Ku7+IBe8+n48KI18MIKfmST1tUUUxFPAZok843IVTot
0bNKSWMd39LrBSZAT1LQCM4xfFw7nDyTJbyZmlJfU3CUrhK1YMaclae6yyPPAEgPd4oqYNpH7VI/
37sC7x6UkGc5dw14iucuA2x+uXxVX16obt58hYfsBbrfEqZGvAS9ouhnAeoRHE4WfAD3YuasmLtX
tnekdRLS8ijrjjtImliaBejY6JGAf3F5ZRwz3Q/eAKmAJ2Ki7jBv0lhdJ5Pyge2GQF3IjpGmdhmI
2rGq9iJ6H5nD0uiSKPePCMUrWOL49QJ6kkuoMkKu2IwHbqYweNmL0+7VXkgdEO71fQpYEZ9MNgan
nUcLFuCjzn63p7xawRhEC0uEH7zwfG9stsR3nKr5pumH4NBvQtqJqMeUIGkiPFq1ISrCarXxjY/O
01bEMTIDV5JqPc6wtTMrDsv3/titvarXRUadWk1+wi4AJ9IS3VtTbNoYTMWecp7OND0TJzeSnICD
sY54HK9trrcWLH+4Wi97dYWsH08RivZzSac0Pt4SadA7NQ7AR1G50LinhaTTmgy7yjdhYpj0dv+0
74nCIEqbQ0Zy6C8EvL+OYaB5yG6PN9fyntaC5LZlZ+SMxtaLuZ61lAKQtEnDUp5sp6FPOHcRsZYT
mah9R3lA9UO4s43MzyQgYgQM6SUeaJ6KegPKzi3z5WaJo+uQ+U+zKguQ8oGYk8vHHqLNaXKdiJWi
IwlfiAFiDCVi/yfeFJZ9HpDb/qk05oLewWCyKu1uO++oTo4142an/758iIgDA5X3etWpXmgcNFAA
Va6IZjdEZkDT7LVq5acdpxTXGpqmloN9Tn9YZdhchRrtGsPI8bv6T8kYfIOveMxkbeTA08i9E1Mf
CntVXpZikvfh4SxTSAhy9aCLmRMyzaLNsBpGMpuM9USVDhPPBiBJhCH3YWuUcSxf23RvspSY2vlM
qMNWSWg8H6SObL5795rkRhcv4XSDkpvK3X6Az91L6owJ1T8TxUP7d5j7ImZIRZWO4KsjhIaeovsC
cWHvERLFj+pX8WEUxvGtwAQgJ8+3iRAigEtK9I8Z4Ua+YctgI31T6qbSQt2bb9ySL98Ay4Usvii8
PuC+AtQLZJTdtC4VU3cZRFBvvoCqg1helMEx1phie6hw2HoCIUfw14DnST3Zd5HZHumMNk+blAmB
Y7P5YpBGJQIMDqHqvEfm9h2XCZ/+2K8Og8ddWu8Gmws84Bp3J6X5NNLub95sWi09lldIYe9KjZ87
FHal9ceMG3rw7j3jB0SyYFhm1s3feTcNkESePh87sr5QkhLJjQ9t3gJBxKS7T6M9NrhC/nM1LvBX
jvJXr0L/62YhodAFrAn2HdNPOGbHv1v/TZ5md1q9yzHsYmwt+tTbNv9puQLYjj7aPEodimzjEpEP
IPwIHsPcwxM7BY9Aiym5l2GdwnduQ6Ly0BNUJA0w6/4WCc6fMvHApLgMRHVJWv1HP3QMaThgO7p0
dcupYm+B0mhx4vemIPVrNXLaeRPN472F42m5I0sDHFtE3X9zc+cWx/JZHCiwMsAbuAUWioZFSyhu
YNj0NbdHQzdzcGYikVxEBfGRCuF68LldIBwFW4P7ZP/xvF8fCs5WF7mI9MZBqDhuc4Ftp9eJHV3E
3Lh2VyZPV7pRKqjwgs0ixZNjT63moYapxTY/sNftwYbkcYiYn0u/p9llSWAqe3NHBRGD+0NRliGS
lnhUXFj5yIzjmJ/3AqdFddvSnD0FXXmp2PSVrDf67wnuz9Y+erH3SSLJFoM7rEnCEQ7n0J0PUshM
ARW8Dn9YcBr9ibEnsOYLFkn7BzZqgWCtRX7IJshmwaYambdyXC8bzku52CrqY2oxCFjwqKQAqFqf
VZN3aYY5eCFg3hRKPVAXpHZCOvrbZZ3Hf/DnMmrXCCMyT+DL1Vty+0HA8p+zbGwNlGqOIdFDwXU9
GB3J2cA35BHg5hobgAp2iNykT2gD02vgJ1oJ/eC1B1wLsZRDDzaw1H6acRj5hsBthTXf2cmbWPq7
QLgyL6AKvEyIgFCzTeHquuhxVZFfBh5daC2AEPm3OfyMH5TSjnQaOKR4w/IvBelh2eep8E13nPpp
CbzNWbXaMIptIeNmVtDgOFa/i/yUPnP+o/RKlcP+/94M7iNsMDnkPgMvaSYxkK+0aAl5GYWolKk/
GwL/Q6JfQH9oinW6odXp6ujAlLHHK1J6egChsNe46KeO5sETeci5rUkUK3HVd3YVYQl3KZIZuTF5
Z75+9N9XUdRf7qOesOQQeLcIMFzYhYywPDHWS0jSrZV+2jN8JqsgWIaKzkv0L+U7JZA2up36RJcL
Shqj2sD/SeHjnu/Sorgd+GlsC2TyUAOHStOKsT/XjA+kgmn5MY7UuTrfai3FnsVeftgP+Gog050a
/hm3tLu9ScICo9xpKvwgIWnjeo/Qyzr7lm8SpRWZVM1GV5ffRzovEV1PeswOqJtu8TkFr5Reu652
Al+nmuls8RV0ZzxVGCarJbm1A7y9Fw5fAaxX52WGgmE6LpO3s9sh86D7RvUO+EWmt2zdCRbssIsg
2UMzuZQJaVLMbL6Ioj/JOg7zqkbm+CCxdy0YMjjJPoc3voxHev5cw3tK+512XJu9IKWsFunuM4Mk
J7OkEKN2pkKrEySJKuMz3dAHC51wbPnik2IBfbdfmBPUg70jI9Hx/VdzpWAMsxOrNPI/oyQI13S8
WjRl24YVw2x7XvJ7/flAQan2h9iV38h9K1Uv0s3CHgIqybehylVf5CDayq88yHaOB1mXbjwsPv1J
iGx10hDy8EaIoDEuLSc42VXpzVoBXKtpfwnUOzq14pPS3wod3Q2oFNY55/X0dUyjIPuw1iS45mKo
wYws5HVMg7vC0ytL4Fn2NopHnwcK7DrUL8+9m0dkGECj+gSnPJhGLPtcmdbkEbqKiYq4Q+bz+ZmX
P3miegN4LlZtre/D3pNdvoObO4fnGcfoMPQ77W98gqPLpz+vdNuNfq0Q+uQqo6MUTqVFg02U1yI/
1Ro8aGP4B8qPUju3agQ7MC+w2QRIiFOrKBWfTVHf9Ga91DBW8P09sw+yKbwdQFd+NUEflpr82Bjh
Ol12VlksYQ6Gia1/Y51QtzrgDHybx9tsxuWyU4VKKf0yHFbKDZzsnI2arzhfxPiH3BpJjF/GLCls
+zQp6ZIK6fZlo+T9thXM49OUOem30mC3uu8BwvDSb4m0u2KYhTP5hoG2ZNROyhLOK6fomVtu4SAK
Y9OXQ3IbMGMXte8D00lz/JHOzrjZmoWGxt/XSAt6niI/op2m9m9hci4Xe9XyrOq/H0qtMWNHECWE
J1zdFo3aatpcAbSZkhbcLBxPMrSASI2N8rjnSkQPrgkPbw4CGF2hrlSN/e61EjMcUZKXmIam9N7B
X4j9VTNt7NLjnOQKWq5xkNz6xsuSmaM357388sMm89eY5gUED33nlHKSARIk8SP1iV8cK4kKyb+B
SJ+rRTILHaGz1nESKog0ijBTl71fxthhW/rfvcKxqyYb9GjjMXYJgSS+vDZyOLp2G1phY4Nk+wEr
33s7qrnpH6rZMlA08beL35RY8Z9rmCgTxuYTEiZ9FsHYzPbzqX31yCY3Moi45qbkzhyg409tjJ6q
K9S5PNlayUpaeqKEqQ7qsPlpsR7VFksMP6zoedYd7L/hmyNYycwzJly/LW0FZt8NDU+nf9egjceO
uj3JzSkeONOVLSKZFcxn8cB3IlUohZ9KDTFbhT18UDMeTJ5c+kclrQiASuplClAxJCxlW/TQqkSQ
PWN5JnXre0lHH44Bt+aL955GvPblFEKab3IIHl7dDwNEsQqqrE4nGhlE02ArQ74TSDXrES2NeZJt
N+4xMLdA5DjC2qu6flE/G9uT8X8gmI6PAj7gkteC9QZoQCv51yDN79fdsmQUNlVgU+NPyGo+50xF
cmpxlHjabYOcf7Fi8t3xstbN9iRDP4cHbGC/GF96oMHZRXdvUi8k71TzGlf1PdpT3Xz4yPJMPc4x
kLdnOqBX/fWNu87klT1wm8AR8imebQTEhGd8fDcr4YRBqJQkslw83b8kFOkNQc/CZuVaFUc5ySDE
hAsB4k9Sj/l6OO9cKUfWFEiWnuHfthX4KFExXFw5YMTZB++sSOBctko0X/Mmmt7yasMGZ3YIwW4q
6srIx72rU/F1iZSl1gslb6AXIAt6i6H2lrHOWuVgFNOwVYHBqfFUZOGzPLnfddJNwqLGVA6YC15S
z9RijNI7Q3JQHCIP1wip6zZ0if4Imz99sSCK/YOnZd8LVdh/Ef7AEHJDUQuAuGIRZ3XGOu5xkhT5
8P8OWkYqXXq+n1KA2qE+Ul/FQJPCrXZGGamCPVEaMsHDvS4n1IZPoOl1uyAX0A4LkErWoigUeDxP
MTgRxw1dATi90EF4mgfBG7ebrsckQrf6rNrjyeQkcOVlUGHHq2HGUVpzsKcHVoa7Hvd5nn8v6qSn
kjd8nm6cyylkBYtLHeotMaD0RowqN1zj0jGn0Rk/+agXAPAt6Q3UOSklWAjaP7pElhCV/xoan4K1
YT1tGujHybNhwp3jLYJEhEUIc5K01Y2bcHdIoLekWUExbDVBbOaT7KX909rBOcKtaxQPbKG8j+Gn
hBzZ/Lx2/T2PeszyytM2/5QvnlkaM0P7cMcCMvmo663sbaululTjDjqhsQm3KL1JZ8BQiR/Sa81y
y/dgd8gJeO8Jyc6yy/k8LpA8Chpu2+rOEi9UTvUplLRPVL3bxM8YzESRkGUcJcROb2mgu+7L+c5A
KuH41ay/AzgHiriS0bAeq+p2acQcWXqckppVYNwZYhB2VOzkuE4kI+AhONEv9xZRhsKEICGI53gX
yHjedgQZQ75tz7IWMW2K5cswSPEJj2u5jVBnsPicHhX17EertB2moUMSmaAgJu/cZuIHI+9X9+3c
LEwnmns6FnnLhUO+FxMqxs1K9x5rp2GR5yxW3ZnF1u14LzRdKN2byKAbvk4EYOPKHK8UxvTtCurS
V0dFwYnVlpCnQlDSE2z63WKwHFSF0I5+uyKkgTyB2ShkdpR2smADsQYL55xhXebXtUY4jsqGpi18
wQihbiQlBquA0lPrw4EktxKl8AbiUpVqPWr0nkQvX230yzZ5dpcX3OCIvtE5s72LtzckFZFeL/xA
KumVhPA6vY6WoX+JIbDfQoVVX8qOwlgHcxZ+sZvTlhXF3+CgMoUXJ55PxRRfcm+yT/kZPvec6WYX
dPX1A5saM1yEQTS/snO8CFbI9/q8loTXmOFglSf+L22q3nZh4Jys6/2OcJeNKXO7Dqp/kc87JRfo
i4hVFgClagbKihPFKP3bmU8HctLQeoav+lHKh93uC4qDl3oiio1Lms/nlKnTRkmoYk8jHDApQ+Zt
3ZTiIjaecj0v6Jw5/iNIpSr7Aw7hIERHK9wezckwsCsQPgPfuWoE+T45C8bzkwVJjmj8VF18KqC+
zk0cn+efOj3vMtFokRBP9bGnY81GJFr7+Eu7sGR/jg/Xh31m3CnsI71aCLzZa6DcRiK/V9T6XVE3
dWB0IRb8zU2zKazrk09KDeUiBlFMH6zUOKCjDZYjpwF7W7+6E67W77M0zgGCeVvL+tOfgUEHzcEl
wYzLueSAG2OhiFiXYTlWRk0g9bDNIfy5Q40URliEU5mLhUgAYgLmiJ0Xbd0QeY4kXPwwofWOj25k
+nfj4tyMFcO4O8A7mvYNatAMAHHg2zYrROeJcNfAuNl5mUItpgaX+TuKUMJSJSjDAKf1Ar6CbulR
rluJoTTfcqykVdlhEK8j0ecPdUhINhL5wadTBhHn6c5QNBNaygYMcKhscF/iw8E3DFRjj6/bc2tr
aRmJKg7bGxAApWqI2NVk94L4pQV4IiSr3IKnX0hVmtCRdP7mY3GSj2V8P5NjrOyYalkMvNdpuPN9
ikV02jOA2jVuQBqLWSpp9b1eZIg36Y9XhavE8QLIkl5+4y80J9jGTd21OHuvF8Wn7hcUh3F8pqbf
jYXtz558XbOa+ddgaG7bMT0/mOZJmfLQnvKCHyERhfDtHtzCni59cv11LdErlD4AdLmnpPWkIR59
0kIXZv7sc4/imp75BJEqetiNOGdhMw4NIW0T0CRHIl43pDBDYo5USevfqrUPrGSpfOAsn35a5lMS
ipCWhaxCJwmtrNi4vjRd4OgPsWVvAPjG2+Yklc0sheTacOYEiZSmZrfwRBxUNaJxc4PvpMy6z6PJ
KBK2ZXA4WTrJNMs+mpsKp9aOBs5fQp1ale7OdXcE9ABn22nZaqAX7suvx9fCnsz3HWXoZwZGIQO6
OhGCm7nUP4o3ocjBebiUyBu9p2NALMqHiCIuJXyYBAwM6hlsheN9NkAgCWPvS7qtw5EsGAQSxlBw
ufmSfM3SXkC+AN5ttJiyfHWDSWOPEXtxLyvswZj2bY82Zxg2L9kdDbEFUMOXlgDeup5WFuVgRNhF
y+1uvULKn7CS6HnkLGvq+mdWKwLCH6RjBP8UyXeh+JdN+z+oKk94Uq+HqIEbkkOt8getPD/zE7EH
oB4v1/cRjXvydA3Te7W7pDHO4JPzd+an+T9fgXpkXibbLk+JE80esEqQX1B5Smum85vSrvsqsYbv
q9CqTOM8CtBu0GE7BR68+bCl10v5Li7T6w2lQHnxZU0/KQbkw+NFMB6a3u9lXnzy+jNgkOeJkpeX
/7Y+jmCbZPwP/nYL+hsWrwU+t6G8R6/UkTOckWLKFqsJ+5IYGeUWWMhND3sZQu0xCjjAjiGYoa2y
IOdDlx4V2lQpUUpwiYwGNQ4i1r6gt2x/0QK+gxz+ChpjQBoG+DjqqqYJr/8PcU8AWtzO+w57U9mJ
b4n93WHS1b5L1+4sQmuzG0FDmpyMy55lQQ2kt2ObKWUhzh7H5t+gnVyOTvTzmZpW1JTbkOm4PVHg
gB59jou+fPJwy2n/h4tZ1K0V7MIHidOFKJBWflpWwxomnVWUOC8FJOWxI5z6HyoJSkYyc/ZXg3Dj
xTyB79p1dSwYWO0X3gmHgZlnrkzV+dJ5UFU7eizTlQAG+wcjoKOSfABERThCfvRZqpu95EHaJid3
5Olq53OF4BemKrzp8RGajLRF0kMiileMLehS0Mt/FLuHFJceVs9Gnk3F8iUwoLqh2v2GlBGz2qiS
BM+OIRwa9xy2lRGQsOVEALlQJlYEpd1wQCIy/bUE0W3ZuwwhZAHZNbEzLGy4Yr8hW5wB9JgbwPAY
m+16qggkMTiipDKhIUv9LhPuH3m3phFuR54pO3/aLkpwB38tNz4lxCxJyGI2tE5JnHtctx3RggkB
VJCgNHc32VP+JZ9AUGsTvyt+ZXDYnc7B8QjZFxTTzLRux0xRhxU3/stp80ehCjyi9OE/OkwYin1V
F7/C2zRYhOHYZXjVKUMwEWac8qVdWu2g9hKiI8hEL7JmhoCxCCrnN5QXltyxjFM3+FrhG/4B8j7m
OyLAjd/F3VdIDdRFhRZyVpT42oumBhYb3xz4kFjgdxeFOP+73WK3EEFsN4540wBuvwhqEtcwIfZJ
61fbwVbxnZxe8wvYiKM28XoQtmm0TRC+MCWb7hsqqtvdQgIntHVH9MdViEiK3T906GkT9PsYq2vO
1bIwUk9rn3Ywd72643mxl/BX3nNdyJzTh2MI9BuLnLUuWMsOTdGwlot36aOylA6odBjkZJmTiJkN
GUKVxUq1tdhzQDua21q/9bSPzbJyTJGrHVi8FxTK00syfPvNwt+D5J5UY4L5pFQQljpsyxeghSI2
mhlsH5ROZf2HgPr65epx8yvYXK5z9XU9A8xDRK9cDBwqE4Pc9oNLVCnauSPIuf7i+WAY9da1dxvX
H2kL6elBhOfYEXc/HJCU84294KsQERUqlG8ftrU2+TPxOii7rcmd+DjxVJlzZstU5QuMA3oVaW03
H40pV4Ng8lwuJd7W4THIPg4/uOv0Jv8UR7hYdLe4M/gO7D8upQivb7MaImVcmyh2n8kLSqdLfIid
goURi5Zvrx1+fm6od/s7XWmRykF/XIrrjyrFBpXF6F0en8vCQY2iyFElIOQgD0Pn+IF2ErqfAizP
I++kO+0G1Vkn2PfsTUJEIamrOg0wo0WmjLXgu8xpylIE6SeMN7kSb7SdVSFVvJCN2ROsmhEDYO3w
BE01lUbIPuP41E0WbZFPJK82qq7j4xoHlLSTb8q1i3WdFH6GLm0MBAbVOvxI+RtpW8L8sOsTsNVH
uZyJ/S+jwRiSaM1gWFv8Ydhn2zH6i9+AhHfooJAwQYllo/CzgvpbiGOEzGqh/UxF8qTgv7YFkkF+
aH+YAXkJRqLd5SoUTK4RFP78mcoL7xsoeSpNVFxf7kyiR7t0zpZvMx0XwGXN/XW4LD/BjjTai3Yv
dwZtUlHfFK/awFUdkdvq2fHsKcRueyVCMvg8RUB7ZCACndopQ5naAd/pLbI5+pnlvYBO4LsdF31s
9bixhCreF/9thX1fEVX2zX3RzR9E26TZV5UGxVh68yk6GpomnLppT8TodeDHNIiPLFzaZm/WaKx9
9ZYGmsPvsrgUp60jBomCapB+q3VB6Y8x7coEYIXD3PSdXeJ7EZWvlhUuMkGrI+Qj7SOIrfAi0BFA
yaepZWvBseOSkNmHnOVmKtbeIGE0VIRvqG9JcK3UeOn6VLwJRzO5jL5JxMWk6EVkjZHOoSw4uEeG
FCbfXhIQxFxL4c+g2iAniL6Ktl0P5JyxTssw6/uUauOiMy9/Ru4PO+xcVI+WtQxK4y5Kp9trW6rN
r4cr0/eDpPpnytMuWY6Fadzr4cVPdbRw9moOrGJWweF9s3/bgD80Yh/aeTXOMZnvl7TFane5YTjh
I05SUSDfhbN7FFJV/ry+V0/hVlc02ZWyoqvNk5gkXKt/pQSlXEBGt5q9HneNCcX+bVltfrrvX8i1
nelTfvL/qzPKZY0e/TgVSgdvd9ZgPyy4FyTwMY0XrjgqCy0y3HBgy0heuYH6COegs57PMj3QBFMR
Mjwbm6lWQ4FVBEzGkKLNjyLgG+rbKIZBULLKy4oqe6E2tyEOC0OZFrsS+qOBHA92p+fn7vTHL4sX
rKP2Euestw6a5X5ajhG3o2d9+zXOVzXLovXpEXzwBGMz6xMDWVz17Iyv1tFeDQZX3MSMur44moQR
Fm/nmtekmEXQCFXEvTBVCnvJ4gfG0TcOQx4lDcJ6OHrOlkZjzawL/HIRPX0Ywp587A+kFSmadI7v
AxNLlzsbDaRrdVup3acMGAjpTrjyLR9fR4giV+nPFnbcVnfa698pE0lRbDtb7QDT5cRh/9z6DP+f
1viU19p46tJbe0hgsw6qrGXWsHjGod3Oaww1ADHPyZwJjRvMNYjrMTkdUutZHbYR+VAWIGBdNEGJ
Ns5stjeWbXAn/1F/O4kCwYIMseYkM/YCnXnPCcFD3rUOLkjKiL+IyLa44kZkVftjcT+ne72/BYw1
BOV3iuyOoJ8OEtwHC/psDq0ANpacXiD3y96oKXZgUm5PbgQ2ghmLx1IvvNr2CyP5Z7ykCIeF1wpD
u+ki5JPawzYHCXD4iQBWSUdBBC0ASjFcOZBoXqscAVH/pGlXy2gLKFFJqtlK4XZQjqP9dVjsoCz7
kCsf9OLBGZkS9wCfTXXxO2Wks89Ex45Xe48+6nTHcdfvQTWdJq5/qKOE9wgx5JCauABaYjvbIxPC
HqWs5ZYeKwvBXo/v4jLC+pngGvv4WaLx5JA3xnwrzlDT1RhYTz9Lm/HP1JEo7wVzYGtsqMMVL4mf
iLChXD8mkv9HcH4uLbSeGFNdDNO4lNo8f/35K8OzS2Xw7TW+3sa3tGMhU/ys5qWqPIF4D/xwv781
5P6uXCSw5x4k5FiMLp9Hi+sYI8dQK5VhRSzAC586KEHnV2nKPrA331FZ1LhUUbIVoYrtqVNcbJ88
aofl0J89Lv55/VCK35z3wSBmN+OCw7mLm0nm/Xa1eDLhY5aqdpXrX+HXAdS3YPU3CRfq2TovDO63
P063iFQDR3zZMU+2mRadKh80vNuL6E1FUDqZcpKJeDbdyD7hnPfqY5R7bmZ9RMs1hBuPn6iUH7vi
AdT3cBd9eZqHQNe5Ibk/dZANWRyjPU4qBDAXnBr2bYzXkD6G42vpXpPjQF00mHSKB8jd9NlAwrrY
ADOY6jhzciuitksKt9LGyaRZtFql+CdP1pOz1m40q1X4GJO4ZFLLn0tVoth12F2ILu9nKs+w7YPQ
qTsSERbUAtrQ2B9vL0p5k7K9HeVnGLFoY8S3H1iIDcWjV+raNAL0waSLugn88DE+HixHIJ+y+6Ew
msNkBsOgyK2dvjr0rJd/LQs4nvRcPGi4jePZP1Hf+kxBZaioV0unDsouX+wqLJBKywcdxLd/nmgq
i0srwtOc8ZwnMWvGyLJ88WZcF67yhNQbyBdP1jSuKHKlU6G4YiuxGQCvFGQfldnv2ZHgpEtBsK5i
R54iUn6qUOdvKxG1qCqpFoHHlzpC30azHxA3d+NStCOvA2xC8CcDM+aQtfuGQcPKTX9Wej3lucaR
wvzbLQ8qOKuZNovS6A0tKYs0eVmJVp7ujEEgs+18RGetu+bw5dozpoujQ8Zu6b5U69/CSR+ng0Ln
OfrlTlqITknv1FRK1yUMIXk6M9pQt48Ypqm2CY4OKdUa1BvYzn5oGN1ebSsT3eBWBbLw+sHfNZdw
aFysKJyDnoQ71uXuBDhyaI90LW1Uq7gCSUZ2nXBYLiwZdZv8BIbMgUwbX/7i9WuSgZ0q3YaUyhYz
bkW5NBAg3kCic9latzsIVPGHIiRg4z3/8UFYde5AlA0aftIZ1bHmDkAQE4kp/9GjyZEdB+c7d7xL
rNcWVhOQafCxVajDeH3tRo/FC1xOtIJmFYhlb0pioJZ3/BVBgd/IvmwvYSS5NGvhZiWf5q08y4me
Yl7qZ+MihUuSBG7ku/lbf+POzAr63fDw09ZSmKSnfo53nWFXDWT+c4Bv7vVUwwKe6+34hoD18eq4
t3IAmJ0yn5k0AlYdzAz9ftyVYb/K+8YM3pm+qVUvmf1j6UJ4fyugvcSEnMsazpAnTjTmNuaLi4eP
6plrWyn3/k7/m77O4sGKzNeNxq5AHi/tV9kn8K5Y6v+n3wxB3qeqED0gAlcED01XznrXzSNisAFC
br++Sfda6f+ldL77pUr3Hkrye0ATSCi1gDqSifA8HbvqM62c6UhK6pZtquJNDHWfPt7ppZRb6Hx9
6qmLA057CDoqY4WsKZPxXZhwwJqEL+IDs9C5IqEHwszjI8S+iZ0tk17ed1MKpXl+N2GPJ59V56N5
mvVd2dgZfQbnuEQY7XyfAQRu4KhoQz8p4r/tvxl4M3KtTmRKdb4PZVfdJBrPf5/fSnDzjifQtB6h
HpGmHHMCfi2Hgtu6FM8ayDmodaIEd0A8d2rc4+UEhZuLqWYE557TcJQMmssPWl++yqFS+DNro+v/
8CTuRpanHvX08Di0oQXjKj0G2ElYCTfrLWgszKzl7rlSfa4aKyzieOM3z+udeCeswftSPZ62dOib
fSyDyv46Lo6VaIFZcv9M9yGoJkDD9E36pbcgI3GSKBxnsKeLISCxmEn9ukhPRXNpfvisaRZDGRBD
zs4KC7zaxIDfY/6E39865XFge82kehulZ+9FPR4ocC0gw8Ebs6CSCVfc+GqJIaGQtmSxDT5uT2fB
tllBYeI9vJ5yzJ7jQiGOGKO6DOmIZSiFpy7VSoIyFRNDeYuBjXEVLamVMHydHVhn5RBzi5u/QAiv
fpTrSplq2ny5Cl17/F3EyCB/n/lf/uV19EQZUkqoxIFKOj6cOmJOYhU2sqqqGS5mZyLobO5JYAy3
LtwDSZbQ8tbaj2VahAC98LHx6D21lG0aWvpvI3ZH0HZtpxm69CMVZz+1eDzJG7I0Yg8b3BiAURCB
9nrlQebAQklpuAeI/+J7rRR8cJFdyKgmSk3P1T+RJIssJsfapkT7Q/OoC3iUi3n7l0zR5ubBsAGF
xFq6uGD47TexmZS33NTRKzjWK5GWpyaNWJCRALX7Km76IEgakpH7tpyLH3rQpDEGV6DrTp04cYn4
WndfQhs9RYW4xcIikwkzMFiPJw6PBV1YwPQNezNDHR2k9ruw3/itNrneV3f38MhiPzcTWFslizJf
cDCIFgcslBHcTgsrHqw9yCY4mJvsivw5Q5ikcQKXDTqZgM2e/N1VguBON1olETzTOMDSnBKmXAvg
LR4MDatsrc4589/J0iX4Uag1yTRR9Zd7AY+UnQ8xNhfXzQw23tk6i/i0xvOchBDGyA7DzLSFgY/L
XheLlYw0HexDVZfE61VIRhxE+0VGZgnBZbRb1HGprzMNcMUK56Uacgj6K9CbCa8ujFc77wJZkP7H
BUZKiXHtvEMBWl6qLZkTOFcWJFNGHsTbQHdmVq8uHGe18tyZ4VwY5gWs9Z5n7wlzI2J7/8VkM8LK
PzSX3p+nsAvVGTuguTZjnDuQg9oQXtzVYCcfvtJ7ud/0qc2ffmsHe+FQBzhAbio+cDjeWoBiXb+3
2THOp3oPQgYykZ/0AeYcU/l7LW8e05mcpfB5ww6vPKe/Ph22dgLtlxhEmCwmLAZQWYWd0a6DcaTt
d7nskMaT0Myu/BpdXuD75z6OMmjKP8jkiLDaIMukdrEDQRrjdiVPjw6MsYe/dw26UgCx7E9jG5Bv
kNp7AYEykYX1YhP7iy1DO5BGHZ+vXtbYm31Z+HFg/9raZxio5/AC45228Eazi3710s/Ir8iIl4vx
HTAFeqYv7+iGpBd33qx1pJCvGH4bqe0ABODdGgqCJbjz2/Efd1AFGBxffHk0rJxd3ftR8a5BEbTQ
TltYqRrEZfTmax0QhNQTrHqc8jBaqvSRkq6b+QtevwcIckhyjho53bO1YnlquYaLIQ1ZjySI4v7Q
EhJAytq6/Uhqb5DdYe0Wq+4ZEizuX4+zCfEB7TjcvGW2utcaiIlx6UXYErxn+TDs9ex7h5gXB559
AEwLpp/f2O15aMS08WneWMrqhCoCeXYaCetkWK0/RMOK/+uZrD/GPrnsOlYt+L5yQxzumh6RhoZe
Qlw+SUS04BZhXYo7Fv+1coJC1K5rMU5AZlECf8B4dwCHiQxyPcwXzvkwdgHBzuZQSm7TLR6wCdJS
VRKzB/ookZimWXNXlrHAulXqU9VmtJDdmEicIdVJ21S8jbRn1TALHU+lPBiyBnsxUl2L0fZ4PFeD
T0ScVs6Kq/t0mVO6O8zm63wFyA0Q12Pa+0U2vjjP8eGk2cnRYSF7xak8Y6orE/jFXbBf068HZ3il
2rsFJ3lA6kTbyWvnjdHnY5vTUo1JjlkWokBvXep1IBYvSJWCQzE1vKw5Srf68djZrD8cANC6hYyV
UU+cXJJSNp+dEZH1Aa9SqWuPJNogJcYBfSqXXS1jO7oFkPgVHfLStjXPqO8V7h4BpvBif33S0jOL
655mPDko3Ex7lmVFwEcDE2HwzBKWyd/8peuil/nOs3wZn4szc4yIM2Ss3DU50x00B6WKlA5Jk1qm
hFcfH0Yqze8ZqzNS/XwLw0FDi2xPKMapoCrvUneR1Ayhy2lXoagKQS2r5Jb1508j3c4uRz0zR6y1
cGul9D+0SiNUAkbmNIQeLdsFDZvsvWI7ppBn3rcPXNlTmtlqz1bvRWSs8PuvRNW8CTxZshdoEJnF
DiOpFlX/YO3S6ZWQulfjV1Na/1e+WX3TumYjBl5/zc6BxfwdgKSLtNRgsH2+wT2vFs5c/OvdpTSv
W3WmX5P9EXwmELBJci3FsNZzZ2ZDYTXM3+cVDVOazDg/9o92lLj/QQr1161kLRthBh0G/DRtmIf/
LZZY4Y7pXNqpmYb7GW5EgJv7gU8gyNc+vR+qUz/Kuf97U2nyNpmS7Z56dy60TU7kFB5sB9r8Rd8x
THpFWe7EIeb3mUw0alRziKN02lxpjZAAmWZSkcya3ZWJb/QqbzaIoZE3T2dcEepiglO7kwMP/MNb
EHHBuEsK3Vy4CqGZOw72+eGoemsHscd2GEWlf6AnnBaROaPgibX9ITTylqr/6acdMVXhR22yOVNI
4EZopDcYJaovwUqGU+IbcSlf0TmQoeUJ4w+uVZFlvEJIr0Jogd8j6C5dKQcK1e3V04HakcLorEa0
6Y7sZoke2rBg3fTe1zRVcK4cD8DtoQWokSLtcT2ZWciFBj2U3b+a3KcMpS30KqFj6MKHRb1vQvO+
9B3JvAFy3kkWt6pQ9DwbAHhmoTtocSVVT93dYH8dFz/CANAsTwChHp/2gu6hAOLvT4PyGcu2DK4S
dBmsfRSsBXduTfkoGLa94mnpqu8RvBe0X/V+g+HP6vRMwdKmGS/v2eRovsV+W5f1+KX/GJBHMaAD
XPnCd+AU6MrCLouNnOIxbsAHJ+8z6v3Xtu3WAk7hEJaf62lIFDpoHfxrC5YQXWvNWUvg+lzzS56P
7GT5fS9fCvW0gB3bk5Cq8LrT2SXqbR51KcjmTf0E44hcKouqx4pu7Jb6c+pk9zukALQ6C8kGOW21
pQbp0EmoWs0OYD3K4gpltIc2KZVjM5BGpb4BCw3mMusdcFfutyH1u8/CO9O2eAaD63KHColVdTIb
CTXZAcwf8N3MquV9NHoiOkJa+fXJUmHVIDkP1UVyz8IUNCA4RBGaiTO/jq8oZr2Q5AV6Ap/zlRTj
lEAYfOg4b07Kr72cT2bUpRCpeDHYXbeBV5FubXP1xzyaHWZosRmdSm1kkapvEbZsVeN5u94BCdc+
/92NHO/CWUuV9ML1JjyV5bVRwSzqfnb6eKDCtbhxqX6Pyac2LLI9DR7rzoFYH8ucAn9P1LfnIYbQ
8ICiruIu201ifIYI3DENQLTRfhY1vuGePr68FJU2w5tYNV+HHFEnKAfqsoXXtd5vTSmYdcul851k
Vru7iQ/H0kEN86+0zzBgy4jv2YfJEk47Ojb7JKK2uqkICcr8cIzmF/k/A9QaHTX1X7/A4LAL6dXu
mYsC4OXjsHqaFRUO2jApqc6pjUrRXlVwJ5nfuJyW6G6snyYgZQA06+Cu4bonvscdvea2cuzh+fgV
RqXYJdZpelU33xGgrQzwZGV/En6oKMjvDpX4rs49MPytGLDiCORK3DA1GSgJX0Yv5meVZMapPFQB
ppjFzXMa29abPHb4Lo8LLJEGeRr94KJ69ERMdGe9hgiDdQh1POjDTF3pRBKys+El9EpCn6CMazpX
WJyFwdZuR/hscBuqG9k0T7iPeAe7X/mrUwjSAXG36kBc7HuvGnLoxsIQYgyNn+qft8g/hauyHHH8
bwHqsam6IYB87gGwvHkQ8ZD+exzZITBxyUGNBdx8+teFdHSaoW3hbOVBiN8la55bK4w3yHcGIzxL
rKiV0GiIcTwzI1dkMEy6zArVQW27W/fFz/vDVBXNCg0AYm5DMoX7qPgajitcnN6z/ljuAl726BFY
u4wE9jsWc/NDcYOlE+AweUO5JcON2N1SH0ShdVbBeTgWPDc/Ymtukg2XAd8Q7ILl4hbSKS9qnZSe
8gmY0Z4rLzYwh8AQirJqLbjugJ/MsQbARTJndXmrxhUzrBuWknQmbHjlCbHEBTuPmja+mTwXHtFA
vsRyYnlgHGRBJoQQz0kBYt3nosBm8iHOWoeuz3Jjkop4hdXv8vcAXrWoY8uOLTM2/6G17gVknQsu
iqDTtxux3tp7bubwhccV9sd5Oe+P3Hl0AdLFAeu4PNjYN8Ppi+AM6KC7zMk+oagkm0CHVFRn60jt
IZeXLB3LDZN+CwYvUNpq/FmufljoI0qIm8Kg1AGOQmhSZYp4T8/QtH/Jbd4bIqYa1HUYyuElDhC2
I0/Smyeo8QONdDGt3vGLpFKnKflD3KX3d0lcflCZ3CMKB3IPlFehA4RZHF2Qglk1rkE4BCIUpLaT
vlnYYjfa+xpfM04S4SFlnoyR29eEpmunPp22Qnlt+WNkJ/Xh6HTm8fvow/rd2G7ZCya+vh8h/WUu
5pn9dFcLREn/f4QUJq1fcxdqy1hsxTBh4z/Jali+NGBkfVHvnB5PiJyJOGGJ43aSVFimIUx26tJC
rKkeHABczpLpOWiylg6ljGHs3mPWh3XukheCY5M4oAtMycqPNWoQWRifov3iW9iSTR0KU7HjU78M
fYwTjLEIKKltuES3xszmAwLnk5H1wiDC637dDQmqxTpcql1ADl6+NtyEsJD+yn996gPCQdwTehCM
9o6khL6/ZzkKg68vL4Dg6YJrTt+T39P/T7+CzDILHemtW0QSmK8RJFWrYnoHceiC9C/rVIhLA1Zw
QO7Oqy9t+2UKGJoxqYOQ7JhBOF9jkPUjbmmUNfZfZVL0/uPYs46KiBlXw2M5ASLhtbqQnU6uM/ql
k1Xy9DBRrJDx24hB4CLO5qtX6qTPMZjFq1JsSs6Bi+M7MCdd01sPLSH2DWymx7YOcjHpvUQh8G4O
SQfgRgFp7+ACgY0s7+rIAJdZ3q58dy4vPaCmg6RWrkQCYwqqDIQZFUZ1JBgPNsB8jy7slhl1NgpE
YPGntiTGugMIrVflXvkJxWgYlyzI1pOg8ZL+fJdwRhQ0hJ93HL2niEQf8zta52E/vYmcUFVsMfl1
a5dm2TwIkgL8Mb3/V85fsd9gNLIUgKzUj9ZyKSpViGxlovlHfeM2NIAFbgMg0pdrEOfqaDTqB+xi
TyZnNSrrSy463zWIZncuIJGhj5wSkU8HoAw+ato2tCKcJgroiFbdJoz7g4rDrPYeKOUlRPEqA4di
wDogaVyBw2+7fnfmJ0RKKt9ADQTEHJEkvC1b0EsfObuF3eTf3p51sQXUUzGUzftXINX7EtypLDl4
uUh0aARp1o+qWflCXDWIDBpS2R83d+ffVXByWKcGdlAs3lII8TKRjhoo3emVwXazIxdsWj1agGu/
Gkw1bDHxNDnAmK6wfv9FZTlI1dQd4vm1lyj3tpX9DTxq0X+GOwlhvuNZGses3WYovDTNk8ztSG1k
JaIOqlPgWstspNGcxZcVIKYE7K61aToW9P+5ZhWfWiKFERHdhqRg/vhgFH7vwYoFkOyu+WrohYAU
xs+5UcYHc0361Psris09ekkt84wdnM+hl1MhjEAsj2OhZdNP0s74OBdXVPZGu3/T595tf4MxyYfU
plc25Vuke3OpBaEcgCDJX4vAitGROKi3Yv89fP25bcGdkLgDvSV6RmglmzPUtosDBzh/fkviuqqS
5XXkD1HLcqlia5K7naN8oD3AzqNj5UhdnMGM5dNwRgYd2Scy75dqLe1WnT9bjm3lrqVd3RhDViZS
7KppzB2bHJUuwL3CInRSsA8lVcweZiFbVL8F4ZugEpWShWOs/UCR1ofRc+JkRJngGIijtMoNc+8s
IdNU/CW2Hkq+JnOXjMWybSP3XXpJpVwH8Az1TJXgZ2Ye5RdOdwfbBO2i7RnJAleNOXE3gvopjye1
IJQsDHTWA+5UAOB76QayIYROW+/qyKjwYoCo7jHqp4rrPoTwyn83JEfY+7UDQkos+CF72Db1lFIn
fF7PLdcMuqMVwNzfwL1eETXfPRGPfoeiOQL1oihfMrTW3leSK9EVIaFQOyaof2qGEAnlO2Z+zU03
aeGMAIB39woqZaj7idDnj1vDNFqx+x6Z7xPlIIwdhYXazrBd+eUoRathcTD5RT3oPHn49CR5cz7u
qj/twmBmi+a92E9uJAFP6x6MnvDCfFcocChxdsVhmiJKWujxHAw4TFe/zsNJ7xfAMq6jZLfQoVk9
PS8UVMCIceiDGdijgOEUZHbbiesuVQsfmnJbepJm5av9jqphh+z6giIUN1gY4ZD/KU6sHIP0lUoE
HJWbzuOZuZCITGwmCZoxpkEjowXhggeZEXB3U2hXVWJhdUPNl8YKCvYy/qojh6MCE/WcUMS+hg/h
IimygGaFYSUO0tIrSm5ZH2xaOBCQ67Gssk4tkwTNOYyyw6ZAsCqAt7dbka1ZPzVzHKDyd3Qiv5ZD
LDptHl9j0vsSI3D7b24GUT+z5lVCMwKFhef5ncpl5+sjBHT4kJlyDYDEmzZjBa5L96njnpa007qr
eO3gwhE1bELxroAugaIdFHpYMooCkPZcyQCtY4XgUIwi4599VLPamUblfr8W4KWyLZoGOtyCKMBA
ezcilggksAUJ0+sFFGFxc7dKnUSYIiCzHiSUY0r3lPV57DnllbUlVMjjiTVIvqFOxEYTqLRTxqsn
mT5Nu8RYnI2hhVngAQUgmAU160hTHtoiLLTEEUSgZxjCeoZqFbk1WymyD1yyYbcDG5/fOmKCtlOl
DYIY1jzs4VYW/+NuLSzzauOyDowbq6vu/JQnYfv3UbD8k0B/9SUleRKmnJQ9OkWn6EjzjGHtGItV
J+HVqcMtezMishSnos1/PeyaJ7oSpQUhFGfSFpvBx3M+nlM8aANf1mL14Z6/4ktTOCkDKcbKlflC
r+HKC7dbNK/gs+c7NS2V1y3bSkAPgnQvIbeA+qVl5PWFmkrtuPZHBD0tDCciTcvc0U6SALXLIxl1
Vjw+uqsM6qeuHuI1K88w03IYxrdE68D3NDMgPYoxEIeMzH0cw01c4OCDZuHnesgZ4xwsa0ifWwEA
bAZXmkCsU/O9S+ureStZJErMGdzVdDl+E2Xf3a/RuwnoDSofJ1lxHko1FiAF7O59A8ODM2uA0lmR
9vCc+izWjDzweMXHxtK/XosnKRRsJeorkFuPCdNBbfp2qdww7SCHEBcTZMtwPhqApyrlR1LD2iyX
EIP3fe6dNZRtIWGBN6OPltL1fT10dCN7n28Vv2PU06Hu+Q7n+ObMjy8KbJndmrAVPsaPV9O5jCfO
fM6Tm0pLQMvaU/5wQl1sG9YPnq4Pmg21YdBJVUzQolVN2ZZc4OGLTPSV7mZNnIQo91VQdV3f7OM7
pyBr1ZKCP9ZvocUQb6j7JjNJaSJUAC/jQj1zF63LYUxqyW3yB5YysfHoVUOExmwZG2d8zAB4FkgO
jLjqeRcKDRG3AO2BxYREaNe6+iA38/Q/GySGgBxrf9UypxXIoOavTlL/Z2QcL+tYG9wZl2Kbl/1h
2AVnxbKA44z6WQiQWz40/q+k8W3pYoROmZ5a9E2S3z5GmEo8ROJoVoJYsl7Iyl0hHRU2Hb5+meid
q5eErgbFkMrNs/m2gU/KZJeQhhsvCgl5xNCNJL0ZuI2klsBqjvYfXtnaYYKH5o32AXsHCuU5WHhn
mAg7TKqsVYyW3st0Ys92VfVSBEPoiobNSS8ku+lyKyK/3GNRqoQVML4IAlSt5dTVMROvXmk72/Oj
xNLX61aooB/nOzJ5L9xYL6i06lpGvbXebn2sOa70QqM4isz1xoNMwKHgZ23mi9mY+G8zxAjOiOV3
DOkQUEzKI0AQbHU42a4u/2VsvAfgbbK+IwZtHNnj8KcyO18yANAPcgLa87fzC8VKsPJN8HMFmBwB
Jfs01hfYuS7h/LXEyrHDfs1oFbxmM2LzB5QmmK647DTRaQkjv0DYAMSrBdqHyw3ubsiaM/m6uqcb
xUX2iOz4lSiMUH10owR7P3WvwM3GBlQnAz2yzuce8pFj1wbdxyovffj+SmbBi3EMF8sQrrgTn9AG
P8macBZUQifjlQocna3ocRGXS4ORPyGpztb8wYrQmIzgVmQG9oAalxv1p/8Rum63fhWbPMBfGFBL
n2aBKtSZdXrd5OexZsm3YxvJosnGAa2pLwrOqJKJ9x26khfx15RMgb6bEiNd8SaD5nqOPl+cETal
f4PBrm+qpr3eRntadZBKXdT4zZgo+xHKD2VongUWC7iRlG61k4+VMngpn9Ft+5FKixZHK9dRvg25
SYjDXws9DQ6LVDMJiITwoyb8Ifj5p0FKAFy7gsP1ZBcltJsiOWRZC0pqoEPSWek0Sd1265Cj2mWi
+p3aHsr8MCZZ/pENRFXt1J0lCDDowLbxkX8bAfIphXr/ICpt28pdFaTO9a17Uc+j/IRF+g/OlfAt
/XoAmdbXRwD2/ozaGHSzyLWKDVuclfs8DzkLYPMZg979uWqAonpGVG1pK+wFw5NZMo7s30/c1raH
kDu7l8JiEfybRmIR27QOMI/Kg8ew//OnfThR/fgzZc+fmMIh0ivq8wORnZw4IsKIv/a3pvwvibfD
kaUl6ffhgpCXsT43gQuYzUqKHIJtzngUhORF2tckTyinbwpAzA/K1IiaQt+My7aWemFI/U+KJACX
YppaZcBXu9GKP7GPVBHPQEl0Zm1wTdhGc3KgcF9wN2WfJCQOgNFX7Mb2otj+RK3ogQvkWCjwMYbT
G/kvljMgVTMYnsjFhWffV2nrDnQmt1knarz/wMjVEWUTTvrNYCGmU/w06U2/x9fkynYhAP0K/u+B
mK7vcJeScZHz/1xJEZeT/DkR0RD/isjhR4ofqtWQabyFPdhc+Putydvd39qErk9wp8fdXPdpLNSE
a5omCULRDRo2MZdAWKwQYiSrdlN3250KVkn0CzqnJvoN1StwWAy+Ha8Tj0SOiwilUgibQWvJVmqg
C/FRBVrKpzBAETQScziVVLivLSvRuZV6QHtB3fcOALFDh5e4Skk15QlfsT8ZyUJqTGSMjruWc9b6
ZlniAsyfIPubDO0pfQNm9XUcXLPJYaVN0izK9kw5wy4gj21O2vou0jIwi835IT6Mz+wfMVMpRLX7
55BIeCvrMcdjkGm7OmwSzUZbCcOP8aTPChAASpHIkjd/rghRVZNx02ApP8KP9uOzx321DyjS4X4u
JoghlOc5uSWHrhB4Gr9C2jZu6tSg1U98Az1fFviioXGcEvJmdO6fbc3G9QFsNGiXBkNSDh1NkOb6
+fOzpRvEemlEOzGYM1U/8dkNd/a6L3eG2b/eeRFx4Hy8Y50EIividhm1NSkgseabi0BrrSl1mfqU
D0vJuzwKZwV66B0sBOxFYzBi9QQSan25663FBtL/uVw1tKiXi/XTIw4OVRW2wwIC1RDzDgP60Tm+
wXGoZbVOUUjJbZA6Rev6RL5CxmpGcUtjzCHcrmH1qjw42Kz+WHca1JFGjRV6s/Y5rVU5xi2dEHbn
GZDpB7pWrNc5UftebSjME1ZNPt1clCUKuiX4iHGPekFC49A5KSoCxolxktazji6g3/0+E/C5LHDq
jpTqW1nErxZRO78P4k95SNndLzs2zT51RzN1oC8/XrjNGR26IfmgBz/uOV+BXdbosy917AofCm4p
E4oHBkpUvGmjZ6b1/vFel47dS1/N431xkZf3LL+BhwjYtQb9bdAm0fdz3bKBfAXyMPt3jwm05Sgb
Dcb4o7S11gbpLLxkWY006ssqxFCVCyfgS1OoqcTx0WOHd4dI6UGbxPacn2d5eXWwWDDYxgLOa4+A
4BkmGiaxhsVJhRFjI4GcXinHTXBOu6vLHaSekNH03jFL9OjoXTPOlGADS9QLFu659zIf8n2LUejd
Jdn2jzk0olC7evqkXIHzmzvEhsPFn9xji2WiOBEcvBEtWF81g93qyT7i0G6Wo+3L/dWDLdh05UIL
2R91++xVznWsSCacSmaHqz+tNpvuEOQslvGZ7c6um/VSdjh+qcKpD43f2KUidl0biIT45CC+zupL
b9xYmxCNsrgkEhQWgcK1UM7i8LLKGHS6fU0DzKhrCt7poKVeT/2V0X6w74dno6UvV+SmlesJP/DD
Az50vK88nzzAnAlXZp3dpZWS6c2mvh4fRqDrAjzHsRDSW+GAA4ejWo7ZtSe9eKpwX15be/ShPIEi
G2rwg9vWpmja655iV/QQ10m8rOlBEjOBvTg6EYzW1CDxucFl7wpAFDkCAj9MJhegXzIIfL2B0ulT
+3Ky7g5nv/LIR+cPQGs1DcNBli3C51WnVWHa22laCXF67DOJn5Sv+thPbTBfWGJw4+PbnvDJs46i
5WgmGpV2E2fz7ed5YbIg+0a4E4dMY0B3ty3V5Y0+rdek9NywRjSr7Sqk59kSSesZEqO2+XaZgijA
Se/z+3HnsbNPCEjTgW6vVf0otukOTXEBdNGRCOigpdngCAf/B7aIRMy7SjPqrtVrfexgCTsUWBUv
+BK2X3UX2s8CWqLocEiBkhjbWcCoIN0uFu7xx53SLBWDDTSRdMex5YGhTz1pb4jM+GejwhO8nIw2
G/7OOZs6u+rs8HgHirkPbgZnO61wABdvUOQKnznbnKPcB8QpC+7j72w+zDvoMWreOO5IHMg+/APm
SU0ykPNrpdcS4DFZdYt7qFCNj49UjpYEHozLZUW9yUz33LKygN1/DZnaPE13ZSG8MNB0Wg+IVoTo
/A1Pcx4mNHFHhUwFiup4gAKGWjmDF3l7Rn7By61lJJFzTwIJQJtPUJaruyzc+speVU1gB1Yc4FMK
3SOGNh6ItX11bijRozY/LVuMZcRqmaF/zyiR8/KHfymjW0/eL46Cu4Am9bCAi6oiEzS4nFNeMWT4
e0LFL4ekwHoK14i6GXqKdg8tJEZdPivOS2/uR6FFLrD1XwpEAZbeQCnMRULcspsNfr8fq08kjB17
AjAWTCAxP4JGBCnIIySEntG4RmJUyZsohhfgAZ8yxMQ7WCQ3RuuulPwfhLhOrnvKB0jVCxBPSOJo
4nfGZqs0B+MuagN4czur2tJaCUwwi2pgT863JErhYE88D91Zt6MrBXVbcYRT07xGT0UM0W9FBfvq
q7gUwtCpNw4yLlvB0BHoijkAEZznewe+R1AjQrl2gpnh7HRjeoYSS80dmzNqLyVxWvuq6cl7IRvv
rqbsJu/4zO55brdFJA5R+k8znKL569IBvMrve3nK9chmxOBvQChjuFUZ/Nmr3RComLt6lXNvsf1K
ubm+gzzInZcQm5vh4AxoFL6+sy//O9MsBpvC9yeCF615JNWgW32OP9OdL/Q8xBv0IyvfHad9Ceg3
nCNlmZmVIFp+JkAQe/8wnkl9bjWA2IWCqX4QvcINViog5oNgL1ViCGE+Ffk7ixvMNUyPvT6+inqm
lvh0FDgrCOLFCvNQF4kbhCBTZA8jKnOi01IXCrU3Vr7Rwzc0k7AKfnmYEqN/NkGEwEJNsLyB/GXh
BMXHMph9heIGWs5nf74cY+nZI3EXGR2UPCtkXcCC054dVMcmvsTYM9jCpiTynutmeE288R4zDc9w
oQur4eO3fpjjoPZmoZmm5HPX8y0Z1lNWaekaVhe2y+Z48kXEva8xJkAkqrJmhqtkvWm/cca7YxPG
V6DWWk1G2TQnA/YL5V4VGom9/jQNncfOHNzOWI+97g91OIz3W+wm59joEyXGUvY68uXiV8+TjJQv
Va8NSWZhQvcwphAHOc867IF750/GZwhOmIG1HLI4pgMbjRYTfFS/6/pNoSaR6EITO9Os+j1pHv1q
DO6WhhravzPzxRiMUlGOhWOEY5JMnCgQNbsV5iajHxy++q16p6u5/S94vJt9dpZfFX5em5EvIOic
gNlwCpdQ6gI8ocGWVZzWhZNU/0kpoRv87FGjgs7G/PD9Q9rUftpdHR1xDrrDrZ3bUUsbsT3GSZo2
5wJuVgNCXBUOuiW+loltWJfFrrV9p2eo4ZMJRmZTyvDwcDPYyqkY89z5CY4sI6YSFpfMMBfkLmqO
QhiF6uDmD3EzlhpL6KFv69iBtkhAyw5lLgmB0oM6fCM5Rm7axtakLnh01yQqbQZzQIVm2NolhdpJ
rGe7ibN5qz7aQ759IXRRBy1PxjFfB6WgkLw8CdapJYZpBHzhqq8QwVMEpbeMp5rkzavGAvBjPR29
+UZGRHvOp8Egi5TZe6yPC8AUlALcHfv/k9W94fhYq/b3zb7tkecY+hIcU9DwQAi8ZIV2lfNEFFC6
jOSsFCXNCy8bCi0KZiAWZ39iG6l4pIcorqFklcS12kZYJkxKelN860p6vLWo1+1JxSVPzKmM63Y/
rqD34ChUUnTh4lqvd/ooNXRfWAuRx/l34QlGSoEJrX4g/NRl2tRjdTGAKy4WU7gcaL6aKPdt8vPV
cqnMjKrTKbKq5uCLQO07/moNDW5Euwu+rzo0tW8l4qDVzKr+CvThiAqLXprvB5T0zXqC7Wya6m6Q
7Tegfl08dRgYMsE0DutHgf/wGIEEqvpTa6A4lBeisvR7VU17BJOAcKQS14h8tJ1Odw55Fz2eM8Y1
fwkO5QpxEXSAGE5v430pALJs84LtR6QpocjjL/3WcRaX+3M4i/dCtExhlLnstIKL9bsPaLLmlh8j
QJUFlOB1fRXt3VqAu8kUnQcTGzkYO6WZCd/ujvwQh7A03RFgEHHc9b0wKvGLIUU3giR1eIiGKoFo
pk3qPdcTsHcY1avq0CwRWKhMfT63rCr4m70SrWp+UgpZfNU/EOYO+egDRzkv+MqN3gY1ie5EWHzo
p5I/P261uWluvLMhLq2d1u8vdAanXx9faSBPo9p3axRHjOeF0ElrAB/W46poAUMk3X7TytZ2qo3y
jgF+7xXpXy34hFqFB/CcFJE56akinkMRX8Fcj1zKaPK1RYjV971H+vO5xheKBY0x6XX2LzvLnb9q
ioclSRnIjJp7iKDHQyBL4iYfP1lspFzSDrnCAB8zWJEqZ4nQEYlcD4gb2Jl4nfsgbqhxhzC/zbJK
3Vxj/jNuxfDret1Eik/aAVbo1HNHhPIi3icnyQRqpnEl4Oc27/IFFR3LYeGXyjylG2tOpu+9MZix
3m9HaOWFdu7jnkCbKy8xoBirM6s1qLpcFooLHjbMTblQOA/1aGBB7A5u+eb9NQErkBQ9bkPmhGWs
E0B5EXBd0UINqPmqTvWZL9QNFmzT7o+ZB/OV2OdOowhVrA7tboCeW1niAVzDSjMhjXD0s0ZtfBcW
q7bnDe7yVVqtesQ3hnyf02r8Z6IMsWDDWsZA74gFg/UN0LmzLknRImabfrgE3eWvWVUUbDPSaUUh
jIMYkLXf3gNF2wtbofhNn1iaKPFUQalQaBnaceywP4ieGVvE8L2LE8TkfFxOEhNa6ep02BHmgetp
4zMNwdtw/Q/uejD07dm0dZedmjKZQFHO0uHHAlS7NEfiA2FJTxIteGNesh6p1JXN4A6joNtVeOI0
8XkrjIcIrI01zIaGuV3lpmxf6n+Ks2QFp0FN/mPcdmm1BiXT7kAqNNS+FwDPQSJvgboRjCr9MAXi
dZfU9zXk5McDCxB5U+dEknyeeiNUIYBjF6W9t3rYKMzJQEJBfTvJ4I5DhMQrCbYNlAcbxkKeg/yV
LCQtnc+tEyBOeNtNUSNo8hLK4MmI+bTf3iu9xFKw2Wknir+sRX0xDVOvp5Cr76PTSPK//fAzKcKl
05ImGyiIC1ef7cLuxsmh5b7NEw6VeV39oZhgTCmNVm5ZCKeY4+M1jnyk/cRexU1A5yfjZeC33fu7
cC2bp5QaFN+LGWIFT0EKkU9HeVUSLUNMca7U+UT5rO4r0tTox86+VCU6SJ/wWaCMiblmfNLVKu30
prKEGRoUgEwH0j88DSKmHl5YJHm7fFdyUWdTrfcOupx/Fs108rmIR+gATYLlg/1iSelwwXnmclNK
PJUfnOrTqEJoyYePdguGdqFbwOV3feQc2rvXJXCMLQF4GjoAFKRxhiqz8KFD8SbFFOWFT9pvh2u5
MyuckAbyAhvX+k80scSCH4VcHRHyyyVkD75VFZNyyNccCKCJ66VaTJWROShQRWCna6Urw8dBgjAO
z0Ix7Ola1mUH82LriNonM0FnK3C1UGdCiEMqMqT6SlU1hGrQ1S0y3QQczRmO0XZleLoecHQUaX9n
NTf+OQLgPbQbRa9Fz7CSKYY3FzCNkihfFGWjpM8HbC3kEJditIHPQnF2ProLitg7F2wL02znIZk9
wPsH5LgCqv0A+vy7vy+sZbZu2V30b5FRAiSqvQihv7osSrhwnEZWoikAFHBVGd/6Pi7ZCMtXV2Nc
Xn4FXMGHnGYn/NWQyU22+ro8HDDwyOBRUaA/aza9vH3ew0YVfY1V6O4JyxbAFf17J+vMGdx1kGAC
08rHelKajdCrCQUdz7q48IhxoZzPlrywK+bAf5iva2+0UpOeaESocNuOlL+5edUX7tuFx6xQI6uX
zhd183lTEtBDodXNVotg661GD1HuCfUcJxMBgQrfvWsRnxHQmLNVeHRySp3wLxXIMlxcZzzXkAv3
a3BXj1HvrME1/w/DX0nRAuHJNIMNru1Kqon4jN8tnI3cuOyy1Y5MkCx7cyJfFiCNfrT3a6Dhk1zl
4FU6jfzLRkydbNqD62h3hv4k50EaYfctwxp1oyYwbILlkDtHFLJpdJibE/wGlSbFjEMxgPkgfaVT
eGEh2TZR251K7+FOLZcJW12yCRWzGHnkLqHq7T+HdTwYZCc3IkUknSO8kIgFL6XYqEmpc9Ac3zhU
g4PPKCKHkOLFv7GILKJqrAUMUsv280BETYGb6/P8c778TeuQJdmSgvjxN/i0Yfg1gaNkynGtq5sP
1i04Z+IhcjTHnP73STL+b4Nirs3b0yOnkQeJXrsd60ZMiTtBgoBCnB5PVA3cdE5iyJ+IrILlaiRf
KxyLGfLsItEr3IZMSDR4lYJyJwac9APVeZ9iOyGuonHdMJd/Xz8ehFYFkAoCpEQ80KQf/DQsJARb
S/t2TYra37Ukn8ZXbDx/RUpTFp9Pwmlw0fcvAzQVBLkbYnfvVcoPKHQmpg9QPk7PubtSuY8ckES3
1SQoWOT8SIpAPfx6sGc7NBAZFdc4H/6v0TQMbEQSgwtbneAEEZJys3ro2xPQUeO4myeXp0lUFa5w
wBagVSuvNwUNZvkXLw1MJ1vD8mtMk3k2WW8JoifxOBd1YQxm8qllzQr4UXNDFw2nPNWyg3CMn/4R
4z1CbGuB/gE2G2JxPwj2XOckbf0LNczGb2FHfa/6FO/0OTzc0WwXsL65ba02hxroY5LyIfCaeRZj
tLl1VRXBizOrPiy7OQnmLJ9bPLrh50MXVNB5QbQWt8C0SD0lsc9SqRJ/kGL7AK6SjtL9AwQvU2Y8
U25mlqPXZ30+GwAgtDsLclKJQKhuE6YTbxDy7FXNOygHgXXkXGHX9WMpY/Fa+9BgWNIHpZo/7jci
9kn0TJJDjH7LBYYVO5v46k+PVg2qaUNjOjWU6SGChDIZjXg/bNM8RzdUuHBPY2QN4K6OudMxzOu6
aSi3FeFlSj9PvnH0HtflIti6sSMP8ke1TuM19+23xKXU5Ub79rXSXjaWa7DRYpdMkbfbAS704doh
eU6sllC+L1dkfzYKCrTWqIrr6g4QjqZgqPfJTZipH3EGxN8CwElwqEgKHHAK6Vnertb2zUtAVvSt
GnE/J4mYvewW8UUE2AEgno0AUD8Iu5Ma+CWXk5xuWU8euDR0c4VGNZds7CDrqlGrFemixW1ClINy
nJq1NweiIHMEEx8h+zgGZCtczHIviq/G7/xdK6VkfDqAwaj8CFlf3dpEuVa9SvfTMBf5wVK0DVJA
znd0Qjrb89TDMhYOsHMnQQCriZx2cpGI7Syphmc31+B7qT+VtGzLcaiN0iijqr5JpWEGy3vTjKqo
H89cYq4p+061b8Y/wTeS6j+iY1UzAhAA7+Z8/N2a0VQlPUps6DMN8fLMYgbyvcSlBnfnvqAOzsB1
rsxvNjQViEiiwh0f4e6VU67x7DRtUXTHQIjOi/wG/VPy5/V0zVpTv6pPE3rTe/h+1NfiFsd3iiSx
wsjou+s0+vA/nwtIsUNI/iyh6FVeL+vkV7E70G/ppq2IldBzwkkK1i8XqZYm7Oe9/I1rl6m2pHTs
aXhHnFOpHK+0Ebhs3Sovk8IiibVPGoUgtPMMrCalOer4pwukpbwYvwoC7uS+rpyd9UQINfSDG8R0
1Nx3CsrPpXok9YZIt5hKr+KgowA83mquBCS2pgg/0IWZlNXsvJ8zpgzxz5s0kMGJWV1NaDRpoK9R
/nOP5kOrPbAIX5JgEUaziHPyw0z9MUs410mVlDMYvPKwulwhiOEpfr0hmeBX6Z5w7ZXrrotFv88i
qhc0lkI0vTrdASDRcP5Om469h5cdBAhrb/8+CpFd1IN9y5fD7i4yuWbiu6dGqXXJLszMhPOfQc+Z
oyKgFbBNzNZ+s+BytRYvsvDGbLsCOPcdmZ/YvglwKqOf+hGVy9ukctyq9iRt6sEPQ6BRihkg7O56
F1WAb+RI9RqeRLx2maSY+gxEeTnl2zqymPLuezs+EJsI5MJvUcbYKfoR+/VVvYTdf7WBZ0Cpn5gD
dC63LAZTlUvMtON0OnTRLfYAnFAFMBG2y43Pm/wj1GgttEEw71g4FHLQ2gwp60X95WZAr7nQSrXO
OUklWUcQq/L46+IzroNAJmS/KMI4JS1rvVVAtwIUMRo9mg4yqsNxEO51agNheoKmIuI6/Xd7EYTE
O436EYRSe/DFLC6OPO7Qda+pea9ALGiRq2xfSunjE1a9alK12BOXfB1TpgJOjIBVVzXWVY9duSDC
Ubx9Mvltk81F2KlmRlDk5Ig8/DqhQ+SEDgFCqdxAIee3Ng33k+bhtz1niJYEC96aC3umuW7fVZRu
1SvnkNUT8+OISO89lY/oaXg7HFFi1hhBN3oLX104zstjPEevKFzHcNPOqHoSWNEYV1q+7SmlKpB8
Ou3nGqNMyUawGrvsDgGuZrNV/2+IHdPIRvEFM/H1EaBGWyLc2Uvk5VoqI2h6vPjKj5zE24zD9eST
neBPPNZXWyJ9g+T2NwYWOf0csbT/gBb9AZbw9EYqnSbD8UkRG2hHaet9L3ScMNlHJ/gZo1Kcth3n
fRfxhev2EV1NGvUk8jIZBWyauNHGbT+1OVY1pSE42RsXJ9RqoYwsgesCHGezHmssriXSL1+HtUWE
Yf2W8a4ofbCVa2f57hsfiDGtwLrRL30jSPg8JHS1SmY/yDYPNbuopvnU1Rawu/5eJuGkmZaAVmLt
7ArHYRs5rNSH2SJYeY4KjZJxY7h9S5BtnQe4AU5YpbtBhyTlXU0enp2dTONC5hFYdNjJAUoQTty5
jXfHrargFnOe34Eje1j8G5rmYOfB04zswilFn54czJUN6yFf2BlUJ/D2SDjjhnL6gQjG4QxRSTzf
eUpgwj517fhPUkcxayCdK++GDPw/pZZ56yUSoA0uzjSL8xqN7ZzS/gR+mluAMlCuRAiybn2CGzdT
Y5c2RP7v3UwUQXDAV0ihhAHLb34tzEz4Z9Mt15z4+CuJvbtN15gjPJ+LVMKv4NulyXZDBT2i2w69
E1MmvrK7qdPJAf+A8bqf0eQK1/iwncJ/k+cZtTfqMnGDmRy2vQiohMvzoEJb7qQc9NaLPF/iQX05
lx7E4vQPs+/Xw9i7mEQfgiYhDqegNMlEzKW5TAM5OuyLzZPvNzoV/DDBQXJVw7Yoz+RmNQo+UZ/e
wjJs8CURDGxDJuSR2jLR6t9YeAHLb3cUDb3BRGTg0ESpFywTgNjtQ7CiRfUC2pT4VLTm7VQUZIl2
Fh/70q4UPZP3PuqRQ0ianaYQjKoJrsjD48vg5/2IuMxh6nsIo11P5M3wTShpApvfnt1HC9xQfLPl
9F0hgekCRMkzHfteMvegZoTIR6ir/1Jfqx8BnpfZW+M1vKgZFMTOlwk1Sbj/B/oxQD1RF3/HdmBB
CWNwz95lMcM8A+ADsx4va/Z/jZ633xypHK3N9InAlePU26wSwZXzyJ1zeIVE0EJ4HVfJyAcHE/Vh
0YFDLkKn/S7tMvnADyGR8C1CjbGcQen1yFpZzD8YvFUZ2DxSjHVEuNV+iC204uLRY2rwWmRqxOFA
/G7Ciga7WkBI8t6sNlMMSikMwKHAMmFswV6PeaTcHal5RmGIayOMA/vaFeolguW7u81RG7WbjcOp
aMjgmUhdpfBdjdNyxKRkvaS3Wq9S45NfeEaN4PZ7LhVSd7Id/s1Wdr1Q0csgWrLTocgCshy2TmdB
Gk+6mOhuVm7L+snQYK54s3MvwBBlCTMkWrzX1ZxCagAlfwkx0z0Iw9z7rEDS/ZP7iqsyabmLLygS
9ow4TwC+z7r5QEhW7reU0ZByKNB42KZToDNw7Ts5e08jEjh5fuDXv1GHVyZP/wElhETbJFbkf2XR
PKdhUczG5ypu5ZnjFsNBSNz0n/RmJcKEyLU6MK0higczXq2JbOAX9DsqNSiIoY1l3Ia4opbGLz91
Nny7KA9WtBVeQ2xcDn74YAvFFUlhZcPP2fcSGMf6dHVjDsN8N3oyWnvs64NMMth50PNndozl/PBq
HVqokiLKTouNyr1hpgoTraxsNplB//+xEm3jzvS4IQmSb6Fdo9NANiZOkevS3kE8TUxNdFshEM9/
xo2WZdidtLw+CcZXRxIgTJaFq1igq0qPyevr11EkhPrsqTJfw68Mi30WBWA76EiSzDfgJCx8zcpV
El+SWRvJSHtxoET/nH8kxQLdzq7IcrsFUsX98MwgFD7lDie8orHdFIn8Alt06EZnrZDMMJ60naIe
yVyL3vGuIi97cBMG61kdxbZnZlFau9jiqYK32oBFgZRhsdmz9bPizTgDOxTBKOrYvdEsF9MraGfN
0Q+LFz8iBLtkFMySXPm4yVkFPV2B7oMp1Fn/S3+ck6vLSZTkA++GpEjDJr8zXokPGBWYM9zpKt/J
1aD8RzwLnHdzMsVDjD8NiA0DWnoImDcJ3gdr055klTi7D7qrDKX2i1DgxKqAWpnW6IPUX6EcXwnD
8OaiBdKV2wAk/svoxEuWA5Z1pxR5pFD9mZjsgnPiurRCkqJqwdKSjXOlxu/lFr7kMEQKaSjQAuMZ
KtUlaLgJvrswWjcvT1s+bLteO0c2jJQzMUIKGpaZals450vv++AElJy3h+M86ub6R4crBJUztsjZ
zBBOHU61MrZVffK+NifSBsXYG1QhtSDv6K/SZJdX90QNuYcaef8QT3Eh/gJUgka6r1b8/U91iJgP
mGwwP0aITTmc8qoJYs1zbpe6/0oc+8qicBjrFg0ZLoevEoEEkwZY7SdiO5HubqazEGH/HaXqbvbH
pMG2x697div9CV3BT26ru4L3TO/WW7ybLGXcXtxiQ24DYpfKGCE9RDqtyUUTojLDFlLwD/0DvFeN
Hw5XgQdh3NhxA4eJAnJSRgn77hF1UFccCQPy/qB2RY0PhOz/dboLKedzd5A6+xGvg7PXEfpcNO7x
yox/uOyqw3C+CIVtn/itJg3i9/G43aZMHHMa+W6bLbL2M6+RM48v2LQFu20p9z+Zjg4jpX4Ld6m1
cNM4uCQAIgeokNtn45kLcXd1PzZtOO13u7Q45CfQoqjeRqQ+geBBlgaxB8DrQIFxpvQb1HcqQwLQ
ng5CPio6oUgbzHjQbL4C8po5xVQa9+ojth4W8dldTI0IoW8xY62M/O1hEnSSC7Uax+cxlj/YC8QN
ofzWUsBRUZYCmAppDEci4RWma2b91L1BjZqwwoS7+BZzCtzS1REvOYqL97GQAsccPAkNulmOk2pg
t2hVXCtFb0OSkUOnGfaFfVG5XuI3WO5H5Ilia8xSmT8XMegniza6PJQiF/3F9yzb4zI8QPl54soG
ef2fvdyLv+zXOYKRdEH5lgSWJdnrhTxUKi2CKzzxuSqoYRlNjQsbAgcjZu2rOR2/z+32f6Z9aSHs
SJTr1si4Nc+rqrY+FraaHRwSVcjDhdAPmoazC/GXxTmVKgmtDXiVYsN0OUTll2e7lPZK8A8nGf1r
WYH9QyWNuPY1/o9xVkNTLlYkpRowAocRxgsQ76W2KNVplI6Bc6OEPR63I3pN2u88sv5FbKixMkgz
BCVhAWyBbspSjk2YLCckRcn65vnyNqJ0G+rCS7Nfa8neDiz4URGJkuzHGKLnjSVrJeJwqz9cNOSe
pDYZTCY4nstUvm2iMFuBHp3uNaqV9uw44HWrCggsRhiFdyv8HpdhUcXJ6jyaf5PVB8g+H7C4AEnu
3lvJ9Sk384cG2TivvOIvOR5I5dxRQmoRcGhdzOSK9++s2vWpfoxSJq0DHFwOlre0JwvzoDFjmZVI
y9bKASy+33ZkQ7M1UzQ6xnxISalCPKa7uRHx3dOp1aznZTA+PBWMlGTGyZT7S++NqgYUx1+hwlWb
yVnf//6TGK8ArLuC16LNhTAoFmPdLNLLXBqLTGDFG9+KEFP7etYB8WH260NcEzonIxhtwSVqGenr
Kb8OnrrMrDcZkwvAMUiKR4NkoYszArbTgdgVHvuCxvjVr1YZgX2JyTyRN4+lAVwGpF3Ym/TykZPh
9BvYxLwSBkjiXzjo2X/NgnX1WIClgeYj/rG8LTFiwD7o2niClQA2rt/uTRftpgGYvH5YsNSXMvIB
ZWLb3tVZna1Qz6fXHmV+VfGafL46tMWn7u5yJO0X6Bm+sNHBdPGedQd3yfrCQFGCVMGz3sMUoUEO
ic4OPDZTDFyErW0iR+9W/M8bT36zZMcJWM7+fCBx58dx6G92KGt43wzHiKqsNDLYSJRCLTzPHG4Z
eoSmAEUNyFGEfS+IE63IRwAVWFdQxeU2J2vHjH3U/lgMdFMABq3QdWPnNm6GPonrYYyD2Crjt5mb
EHdfWx9BWM8J8U3p9M/bWQ1zqzlx479sq77Cy6EKH1ALZ9bArcuzVIxV3ESy3ZcUzCggbTTOndP0
9FbVXV648uo1pgNN9zA+eCI+gl3oc1becQsdevVAD+ilfjb7g7LKTVjfQFeKwHW45fVXX6mIpXGm
6GytnBh3iCUTlPcis+dBKMLEGn92obqrQVvUx/n6wu0DXLd3hmDN18yN/2g5MWLsZxcjL3qc+PpQ
LaUFlmqeH2vrsYUxcGWB+/fxF0kDZ4vLUgrX3/S7dFEaGZwDWt2NLXi/XmMtrrOtE8tezS8ouzbB
hrr3jVWZU8BC9xh0NJBtE9fUxBwKa/o23U8N2RHcu5cPPsJ1vq9u8kl5gcXHRlpf/2svPHtPJFZP
0Diy4fQa6H5i47FtzUt/4APF8uqOBWCo0xb7WGQMmy/8oJjc97LaJIg9SPIdYd6PYv3jz5WsgvOx
96nQrryoono5ZGsRN8zGQ1czgPJT96Z8Scjx8Wy6ess12GtjR7EPdESFQR1j7yZpqsqw0V+A9yc5
z5BmTQ+RHrgUptMWMUJ/6IysefPOQLObaBZCeShBJndQsD3s9tahPxVcrlwZ7qj+SXHb8/LVmyol
DSVLi0HBRCxX7rxvyCOOjDleaBRbku45n4b5Y24WoxlyX6716ZRIZf5hskv28CqLLeJqqOf827Gw
U8oG6pOmxzL12SEzM1mN4PDVEQvX8vnaMxxjN9CJXlKsUJt1Bs8xDEx6SrzrlHnn21ap2LW4g6aB
2LZbgsU4nhlgVvIr73/Ditk6XzBgPN/Qoj4bMr8pQcsNikXvsXgbQchduRp/Z1xrDavlZCQLzvr1
1H58abj+kHgtpJo3gCwTHr+ZoaP1CaEbbk5L9b4FlnxG0FU1BvtpOxi1Kr8hX1jJM8yUe1diJs/x
3dYTY8/PoykzpZOOcvEgat0mk5J1712kTew7LyXn2F8oaSV+opY0pnQ2o/X+UuUPloEUD7TRkAPH
qjEzgsbwE4wLLQAh5P2m2gy1C7JLKUCDA12cvGkAw1OLJT8+kYqCehekAOZ6pO4HIE8IzKrn8cip
54wicaXRWcDsbkkKB7YW/xbkaqc9wUxVtlStDMslW6zn7mXOkrgKArWjIW5G1k5vspI0kSbn9iYW
hfOUEj6SmuXcSPJwX7bV0gpFYhqj40aYiTAdZllnsyWKcrgQjzS/LPwHyFuCPayaaTkHnbbYY8mT
GnyO3bHt/2Mx0jwqIIgqDIDXlMWTjDCuPhJr/4gH0ql7KiIQlKB5mMdU+KqIuBscPDhlsMRcH8p2
effKJe+nu2Q21PnKvHM2uryRGAYIiiypE4OXve2rIMfC12s5v02H35hxfMEXj+JrRVwdYOOZU2ay
x46bFSbUksdXOkuPoQ3p/lh2tE3Xbdl0m8OjsFzzqkmlS2AL+WJ+cWsaNqXJkDOhWG+VNOeDoNpx
vJFiLpsZonPumiFa6Zcf6O2Oit0fDReGafegRMyGnJ2Bh/7fUpO7r97E2tchHW3qyk9de6QN7UCO
9obwVMmVwh1WdQCwKyZ3HkjhyPLrWckHPthVF+NMzIGPkIsKZ2IEs33Zw0Gp5XbxEP3RRQz5zH6g
NTLTs6IGfEovhuLReqRrqQrHrWeR4liE5kq2plWs7pg3erzMlGG8nDLPI2Z3nopo+Sb7aKbLX/If
+zCLg2XvScJEVm5uya6JRKcMKgKLQMqNMac7oKgDFbDw/V44TDf65PTVgif45KA+cTzl9C5ebjRh
Ceeec0zrIYBpLPruVHoyRqZfI4qsZlPCaZPpxJVLCap/6CFnanz7SBBwGLbneMVzuNmVULtLhHVy
4DIaHDIJSj6ueJrjJh5OZumM0BT8Dr/kWake1Jb3BXHJ+6pNiPz2iwWKDiFFOGi4/wT9uNj7tVRK
7GxRQeTTGfr67BAbZdkwYw8bjSzyFowFOWye6YYIPSKQiqRHY0HYayJtSiPqeR/z2lFuEaCSHsWO
A/nxzlcZAIjsvR61DgYFlH4gq+9ZhPHHNNkl28NQjh0VHOy8YTMQ0Xvw17TWlRrzU2jv9QbefS2E
YSur+sBdFvJ1UXFspt8gH25UhhrUaB9ld2r8NUSS2HT/8VSkxoVAvAEpvZx90e/H/HqoKNzOzrGQ
PB56XRuhtbnsAmr/a8zPHzMe46qXnc/04/jpMZjYUz4XCnrHmqliYcqlSSSj/3u/TkS+YA2p+HvO
kPf1irb8IiWfJR5otxn8YXJbz4l0OuhBD+cXgE9Ouk2MfgkGFuhKMTb0/wH4PhHkj4CbgbSCOoic
PUJuycGwBiAyLJSAuKySeycauG9pGMOEc/J3dMqWnZnBPlVGS+wJrz0qU593LfIrWXCIyabUz32W
ShpqNQ2yFa6EO6qeUiVEliVrewbGIGvv8PCQoz21nL+KXMqCOmiueWjjzOa3q6hzlMU7shLBYDa6
WJk9qdAsWgsA4yKcuiy0ZYdVjeryb2XrrRRyNqcMZnp+VDGDDcg4tSxJjMVvp9zMI1OOUWrEED7V
IZPRFF99oesbS23taPilMtWlwAYWG2W89QNlBUvf9AiUN+TUWFQPHwNjxgfDvkr3BbAmY+PGgFWl
HlTEcLXzL/ssl6MImsImC3qzEfOiAe6xyIS9V28fKenXiKow3YyyP9JAQwpPvkUj34T4Id06zqtq
bLlZs/unyRJ12nrKRMRvD0F3ms0QAD7BN7xw3qyIyFg261arpzw/mYpODsqDtIL4fjFwrHK7IIa1
VCojqGSOg7HXlXm43ocxHzyoIQUuoN4zpLWVhZfBQUHOtHDo8xfpFgapTR7mo72ZFi62W3GyV6jF
D9oCBiG3hdvZpYFQLX9E0cKg7F5hD6piIQqjWmmxSTiMIsHhYM6qqQmt/GrHK/poBE2Xh8RDmgkW
VeP8KV7oYNb6pzhjb3WygIuGSS6l9XvhfHitjospcmdfrimXN/3qFMNXDqixzLE6eC+oTKWHv3uB
df2sDMHEvJhjlo9ysRAWqAu2iEKQ+NXfjT4n5qB0vo+AK5u/gEJT1r+/N78fS2hy+boebnkiRjJP
uqx2YXqOYC+OMqgqWt62wdr9aqvZqugbMnL8ys7I/ZcqdJ6ZOsOFNf7yAO/Brb8L7o5r9T0z1SGB
FY/bg3j2Ohtgx00IOgnZCQcNyEUb4ya4YVBfUsIpdnriyLP9jklaxUTJQMNOKblCWNkanXZ5dwv4
ABCw9luKbwf5OFwQECd/JKPe+8qypCvaWqbQXlUQnsHfR71QPxbix4d9BwXHMTJQv8FhMJ9RlS1B
jQpQB9TfJr9Mqpg5KYIKvIvy+QEb+XIJnC9r+pQmilCVKMjJCru/C2bwIs/71vSNFVOKULGyDgwE
oTL9xtGxy+Ik3QLeg+tZy+clKZoZJ9bSU77AM+9pZTGnTaLWZvf+S8WDx8+NaDKDTtrXo8OQSBSG
VtEIMmd5Mr6d/OLAACKDdB3O9bC91dEpjU0BBOzZFmoG83Y/JVjN0BkpNsIKpZUUV092pWVgJY3S
vVHydfNh6bvj9EGmGZE1K7cePkZO8roxXs2A34kj4djg28ZZIL/Fn43MygsJCS+dni8f9hcUeQAi
iAfLyjIuBPMNc5hPes3ZajcyJR6/6aeFvqtJgdS3yokNGEs3YaSUQrDfw3RtqzkRYqLU60zDbzKY
FCZ05REKSZcha+igDYMzEt6O+2JjaI1aio+cWgvZF0m2mpsAfvfPsgqFAlYp7Q3jOGnv8bQgE7Nj
IR9PdKvS8hFqBkp8ynSKTXoqfNizYSgtHPELfj8v6e4fKGw4dexHEqdZBhtIlsBbip1VOfYvrqFu
JtaAetmEXnrqpyuwdC9sR0KpWHKHIKR5bOXnDYa8V2jbEEhx0tIHvfPeG4PvVO8oD/CwtlkErgxa
/U4F0lesmOIrIDw2RhzNUmOD9846fF7Mh7snI4WRCZhzKOpEJe7GirAzYOMSVtJSHf4ZSBwZRQFy
Pch2qlO7Zd9SR86h6wangEWvin4nPJHuIkuqGhWKsr2YVMV8RRMv6JukFXtiij0lwzLSJOoN0x9W
CpiPSVlRbqUwd+oUnRAfvy2GFc/CcfMqRaLU/lZNx0ThMt/8a8OsTBL6ZiauAwj263MWRcY1I0xs
UasKITerXqAuGE3XGZPx9Zl7Vp+l5I32cQaOdRMN+WTGaUpyj6bPQbgYBWEIO1wp5arKlTQx/JMa
57F6cFQYaYRBmGnLUiuNc+n0ZevBVnTTN2hllq6nT/OnAO/arSNecI8pVnkx5IC0vsPpE60T5cJe
eHTU1fNv3yBsN4u6lAbTCGYSaW0F4Wywz8tT86dX/l/EL969cSKkFry4IFLfjHRZEvm84v5Ij67E
RcVAMebpqegWZN9+hc6oM9fCoIfRZatstXjyEhIta8XdQV2QASvI+hgwF9NyZYa+JZG1WUnMbtYz
nedwT8XwjNfDpNxAVy7ThG98yZo/mjBCsHYjCw/vlBoPF/2xox7LCiVrHQjTN/OD2a+Z3IYx3wAI
0tiZED3huw/hvoZOMd9PGr/zFW5k5U6KYbGeGhwwf78kePZwxfJnRz0prbW45BLQpVi7eCwZNj93
V3ipAvhy+/1vJwoH+tLIXUU+DCjxEQN6TD1wMlF23caQY9y1S7zCN3RlAAC7t/bEZVDX8046SpBw
KByEh6KRKUtcYaW2w7mF1rYOBltUwBtWWgv/vAeHqJYPsDtukItCStZzy5nUCWxWWfOjY/aeI9kC
dHTI+ypYBWUFORnrlYZFcwI2SEbAVecxjIN4fgZp9v8aAYBQLwZ23OdOSXeYqSQrinEWsHH8H4vV
zPMAqjtOfehGUaxeP4czwyVGUK9MgFB4Gu6RDYyGMFfu6njg9R6Dg+YgX/XOQEMNrDKUsMqF3A1m
bc0bra1n1lK8ZT+nIsvd1QgR7pEIKvSdDyuOoB4s0urkRTdpryUjAZRsNW342Df/iza00HsYcqB1
U4aaZ+keMO/UeMRrCMXsp9DfaDxRp/AYi+Cz5FaF0HrLF+5zuNZoAZ5FnPjq1wzRY6Y+njNOfrGa
PuDLeToga20a2mj3X1WnzveRtCDFExqQxbv8r/fkF9kEbN1XWNrFpH02WkolLTlCT1cZrI8h/Ubk
AM2IPIDHb9W33wGR6elWQFMD5xaPOlp3lIip0+7P8FztAEEndSigEzCAFNAWiYbJWLWiDVJQ2J/q
7Zz2vjqpL5HuH2YTbVA4iWjilz5xFSJbfRwf6eZtjM0xDbQfP4qwcRMJKWdoYgvFvfJFXBzSvhcs
1zjITBRXuNhmi5W+14p3fqEt1NlypPm7xPE8VK6EmuhcgafvCy6HYyl/ouTT6cmm6hayp0OQBM/T
9f/+WFYAGzFWYy6TEwbEb62WmWd/KABag4G9HTLS3uEFgsu/8n+KYtvvuNFioYlGbztUlhOQ87W0
iwbT3G2UBcNQVBzp7HqvEIJplRie+ts0YuGZGxxmLaOYprip2r183UOMaT+lvXJVaQ6fV7texdbS
stfYCcIYcTMmp48Ktf7f+XjuP9z9usxgBLxmkhp1OlAAM7TzksyCnnVlTqVXgn0CqAah4ZWCDtae
CYpipqppyMMnTl2sMAbESvkmdw7T4PsxO3tXsBFkaxoXtaET5NoqnHEeWga0uYTUHU331rR4SlQ2
4/xlLTrGMSg4UBKSTxFrrJ5n7SFVuHGboe3LrUlXaHoOxuRLlApceeaY2wu9quBBWWM+H/SN786Q
ltAWLML2/9PTJFAmQKg3yThtMdjUtQpck13hABBLc33snYFTvbj7whYb3gGjWEfSbbsEaZuwfeK+
CtcqKjUNfKXVFxLEIx+T0phdsOpdmtstMfrjiYai1ez6jxSDYAAbBmDTNIjX+tLFmhMEPFKvo7zx
VcASVTiQkAos1JKwnSxrF/mKPmIBHi8B8EIWl43CEvnLtk0vq1547NB4fudYhFBd4LL1W2fsuVVv
bMPZrQ868eqvWmLs6T13kE2Zep97vFD6ruU+CEgriW6TR4Al4IHzXq34S6oLx8KfC1y5cyQm6gb2
7H5zbfNJRpXNQpvtr+Fx1gYtoSOBTQBSQq1oo9GYBgHduKHC9q8UFTRgS6qq7bXixW3somfaBo5q
+MyVtJXCJpvMHhkkY7BMjvbfdDX/3wAXuTdb2N2i3WZF4R+gIvlkTnK707rbd2mWrJD+u+z7z7cH
ZXFfvmLTfD8Pel9TTT2JsW7ElgLkAbb9Rh2gPCUBWejg0A6C4UdccVz7EbtmajHfm6f8sgpkZ7i8
ElBs2OIsaQ7DJa19mWz/sF9a9zGnz+4TiAJ0L1mR+PW6WJK4b5frYv8XWNwFHvdeJLj+0jz3aeRv
ZVMEv41dahKOvhsN+MPTYK4Qj7qiFpGDgPkvrSKl9k57cvOUUTONR5TFc6g2FCiRr9DCSc+muIE7
BlLxFOauOF0StVzx8Q6mMX7X4y46RpE7giMz8P2cRMrTQ24kyq/WsJylmH5q2Pa1aVS7WTlecpm4
QBs890ZjEBpZRu6ESePUtIoV6V0Pf3M5lnNmgkEIkco9n6p0kh8hR705/t1XCIxunrdUPgBL3PUu
6Y8MCPNammWUgtQijk2hawfKyud6ZqG/d1iO55RUoROyTBh8zPOn7r7qSuHv+mVXtiu3fjSjLFSW
SWehDvlWVIaJRcqkxLIUgs2SnaYh7/I7z8HpVT3WUtD9A+V1EAg84Aish+IEF833flGsQIVPBF9T
9xPC/EFuKIRpiHzFvBSN7D5mDuHUJxEsxcYX98E5c7g4Fjj8rotrnJu0Rkg8GVIqgyd2KRttQYmO
cn6M8ZZTBS8XGY/QdCk8xMML0jyRASe7yTnu6i6EEqEarldFliMziO4OPQXbHwGMKfXRa0nFcwAz
R0pZGXRGX/fWRF6bPcRcmsP4GYwgU/PsZU1feEq0txolpaoAyuFubsnM5F1pytaX+KS2sQKjrcuD
fMbhLOFDrjBxYP7PUXwu4hfNUVn8r+0dayToIUXH1j5A9v6E4J1F/32v6D+nvnj+pgkPbhuvisDz
/cNjhWoDaVLrki0n90BLpXmKZrgCAtth3hyDSag9Gm90pK4IR1PMO8Gm8gijrIgz+q3htLZUiyQI
xBeOwhdAXESgwREun2r5elij/ahHQHBCNazHF89jbRvifH5qEGUM3urLBpoo+hwzNc8OCM0ocKGq
rWBfTRivVv3EApyFxwGufKKHqFFeSt9jRynHIA0K+2asK6jsVFJ2soVr/fZoWuBDd0zsUDMgw32p
XVxjeVcI7PTRQ7E5tk7SlSsENQQkTSWX4dB6Y45MheIidJgi4xekxIo6SwhsfMCxFzJ8PAOmHfIe
x0XA7XPB4wJzW89qmDs9BUycIDziAJFzwJEWjtb6nxjzf80Mj9HBuP1SKHugzY5gbC4s3hEAUASb
BtpUCF+uDtTf/vIo1DTenk8PxltYRMe+El1TtASpMtt1jDz/4fUh2yeNPR6pQBCuQmuYIuB7gx+t
1Tf84JIp1uQY1FJ/FDQTg3eKxjRV/oYzH9fz6HftzmJxfcnZHMtSj00X+EX/G8o8ogyNOL95JFco
FWtdj/+wmPdf2IrQdbhAB3S3/Tsu24nbsOiT6CmAnZ3hKiAS6liUtc6nRVfkbfl2w+98Az98pjnb
IZZDIrdNr42adF1BEBbHYbMKcqD7d1uK6UbtIUUZdbM+fD3Ycm9H51s7AP/PxRRL4phWu8vjkPqW
xf/0erMdG8+mDsw3NZpVfTvpIBmZ9uLgKbi8mk9Dndq0ZbSJKWROPA+fFrCnCIQkcKaxQ/zGL8e+
mBZxgFmjzfqDou6WpCb2ZL36s6dVHCykOUW7J1Ml6N/elkG2AJ6ka1E6rOT4GJqBTp/QmkUdtnFN
3Up3cRVhCVgdc+GU2gvvVKoQqwcJQ07JZDGQK3Kd4gp4PR9cdolNl0X8wbvGMP2UWTs9Cay4+/iq
iPVvk2lbJNY3QnTuB6Oj14ctlLIe9I9IGCIScJM30dHKd745Hw2g/TKs3xyThTajHr1mLnzcLxaY
NoDG7flnfQyrfAHmh1bnJQAoaE7mgCmE4njQrjVqjLni2NgZxBVMJZa0lwD7TQHSfl+GiXmSEhQo
fW8X7OkJrwNBawmr0+5sTWw+0qSl19BFF/rPcKRFJExfqL9pTvND9WOMXCb6Z4Z0EUlt6Rl/e39H
/W9OxtTtokDQrnIe0IfJMD0V7jEh1T+OuT+6oEZyrdlEH5Uzn2WXsx+DCqAr9zVWeIPrW1LnBCnn
EofyhrSrXx5PIwU1LmWIuJ5OucsLn2S+NokBX3faWV6W57oaKkIEcmPxpqz2JC5lVlHnsfHo7X1V
NepqbHaESzb+dharWRCpYzCFNTrS0GROA04I0f2j55BG7sKHRsAgHsl9a58qRFU++/CsQTTTXFls
IzhzL0JI3QvcYNhMdNSCNxQ/U+6WCqccgW/1OYLPZUIBXQmq90yHzUcUPsbkn9XpSxFF4CvcGHfB
9g7XmACkrIHKqiMBAio+mFUN0+RlaS8pVOvQFx7JKPPfQiko5LKi0MJQvmPRr/LEJdYKCvTQFvmT
KOS5FkDDE6z6cmhirszSk84waAHooxRnvKjWOUmYHfAN3DV/jA01hdh+NA6/91voPMgQYhvW5YtN
VCrbRYNR0HJU4P9rL4Dr6bakLy+NlgB5+37TGd6LAa8K9ssWvx8nHvufXNXO9Sy08haaMXTN17RB
Qb/mhJhHzgy2dvd0J3v+cDBqjAPZteLyp+sxWKmvmcpn2QPGr5GZZWc8AKnH6QbJ+8b1HYUZOen9
n2SQPXRzwlhO75ouVMrKmWF/ZHDTO/eB5FpJfk7PA5B2YeumX7oAOCqKWPn9QIN1Qwy6pKqlfvXi
Bx8qe3dKBXfnrJfOkRKrLut/hYNsBDCCi6H0iUp3uhsGVkG+GL8i/8uBVEDC9nFjJLJeHlTeOk1T
V5xHEM61q+Iz5SYgDs2BVVF7VJXD38XaU75aJfDGh8UN7rGmqHAvfh6KzlDsq4f80m1wSKYCkHD0
UJzj9XVr0oavAtXObuTEiA4eC9QEUg6CP1TLzsM/WRrMHtv5S4jt+hljg27+PQ7TZh+J6S408lmb
YXSTfx1zYmwaBE3hAsUmTTHm5gJgYBPyMl04xEUUHQfZ0TPYhCx2Hd/uClzgQBxFtWVtk+xX3akV
iOxyI/3b8FkbSFZeILxeEjkg8T6eb+Q4MuWzUhb7cYwMdMo52ay5lykV1Thl6qS9HJSAphh6sIYS
ox91SDfffxCnvJEL5tApnVdPPn6PwFgo+OM3u4jLyNWAXYOanCZHjVFkrAMPZOKIW3966XyK+2K1
eI0sA9mNafCH2AojWVU/fb7+ULvHJ73/Uz/Yd3F/tZD92SekoygdkH/r0tLGtYuGocjoc3e1YbKM
05HuVc7KW+yznk+IBlmHOwCEaAaNm2D5a9ee6hkD3HU363+KTnaRu6BdaCGcdvubq8TGOyPg9rkI
cJOydLpNRwTG/4fAOzMY4XaSF0kAgvExhbo3aGuA5pmO7p+3riTF2M0ahFKd5e5fYUr/QxGVQ1z9
Db7OqEa0ROTnUDXXbBMioQ7B9XuKROcUOpKc8ScPLgSUp3OMYadvH+aKNL96MSTJ5Xc5pHKAEmry
I7YmxOKdz5NrIgvUYq3drRi5XdZ0uUwDS5ISHibGQglfFOirPCOT3/omVDXtWZU/qS7nH59S++OJ
zHoeKJpd4VugitMy7mmaVVrjzu4pQLhtgs/XmSpaXCTxz8tGmpfZmPwIdY0emakT2aXk1i1QeFzn
EeaJhu+KGEEnVgi+OQp8kqK4Zl9MFaK4BMQedSt+eTGCsrLFvF2gQzShBPNCRYU6ybZm9KdvAgwt
dVI8NzhlY0nBJo0ynhbNzemB9twjGs0g3KXrn6+KsblQbdIYOOVpege9Q17hCb1p21Zz9NbdlG2w
HUpyRLAUd8jhfsxWlbYkf9z75SuYZJzJ4UYMDFB3Sj1gWdOCY6d8xovP+cIinzg1svE2PPqICtzK
jpi78nlCRwBiIEtX4EK3o8oMjV27BagRvuK7pkfZdm8+VR6LWJowM+KpmCCT3NyrsWHfNK18k7/h
VwBo7J64Sum/Y75Hh1QN5+h4/xetCoO/90Nk9s6ZW+TEolV71L1Y2AyQzwdXdsMirvFR1L+EUqDG
vbOBtSHScWYFZO/gTMpBuCHAEb76Yv+l0twIQ3ws2WpL3rK+De6L0eVJqze7MIwkWrOzEUqPQ3Wl
FnopMace4T9GoL22zxY3d4zYHb82y+/y4BpF8jE8310u7pU/Sa8rIrMJyi9E0PRRqapXIYYmmian
HAdCRIocRYl5Sf35t89KH4fdXGojjkFGa4sCtD3Im/KY4LpAfWWfu6wuioLGibFq3FEPbqomRSYT
afT/3N81WxMfTw4pQZPNERqBhaPdh6d9oGPqc7X8u4i2CrlqLGzirRRUHuKXiEf4BuTPcrxwAPd9
iIYGfktNpL6XNi+Sc5iRNSSkKDl1/SIJOj6ZNecQ3bkKoz1+A7QgHmf8ZZTKYH7YxBwmGJmeIDrd
jC36zo/r/UwRNn3xCVMk287I3OMRKmqhkwI9nGX6+Z4NxBkiP3vfDNbMQ/SF2eNzoxhGTSWid9M4
WDV1+trnjdEa1vJlWZDx8WuE1JcCCKsCoKNM558qSGssusx3bfHeMytD8v2Tmd2EbuA689WxG1nn
Nvoqo+KumOAzF9DQGidpkjWNJMe7OENeyiWk1895Pw7mQxy0XHQoFP/NtpCusMkUqYT91pDrZseU
D16/P1Li8toO2uEAC2ejDOdcvhuPwAg0GH93+nLwSuJ28VNZlzZy4dzQHIVIr1TJz5pgnvgeki5s
pa3j4zI9JbVf1fhbYZuSyjZWS6rH2lF4EPc6Fhcp9pN6chwWFJXCwny24y+PG0jmjCb7z8DXiEXH
fDsAC9+3Ydd5d0x6UgXWvMA3QrcEgqSGbbo65N9Z0leOZHKpJxW5I7HjlUx1MmuUxZaIKdxoSDf+
JYBTy73x31afjjRAK7HmKF6tn+uQ/oAQsTxRgfZbsz+557baLZa3tsPQKIxKSQv2WvhZ70HOjYn0
cS6IYQizLe26JhY8KjMvAFA1pGl0l6yHkvAtphGaHgOgN0cXSBPLMKRoc9X9ANVJpAbG8yo9aKC1
CXQqzXGsESWhzthtUB7Lt5frZNDKxfcWGBXlp1flNgDk/KGa1Xli8xetxYAbfPHdPWNJQ/Ub4A4m
MZEoxKjQ7q733F3Hns2WLoagmyXUsUVzgcdDqhrHYr+PCnhYOIQ+q1WVHUTa3zti8on9oAnYIoFJ
KlfSpf56Bvha6wzZQLSalLb4vhY+vLVFzfcbRd8OI5MVbwzsiC54PSo2FZPt8H/VcFm+egludq6W
5D0ojF0WXYGg6Kq68U0C+hO8lW/7aL9dKKnZ2/7GTM9L13dMPTZafo+ZlMdw1w7Xd9QPXWrwqC1w
EObfxlmAZCbx5lwkTIGHwEZ/OGyuJAfpXdGSlcZsz5zvNZlps40uP00ak8Kb44hBR+LecGNgqK7w
+4KWxO+ol96PiS6vXD1IX634y+0XmCiZ1sLVH2w4bJYmlf//gsBvZ+ERNkSun7VtLdEzoi3DCLsr
6SaOnyis1v37fTWRVRl7z/oqdg/iLvaU3Qpashg0WLWSX37FoYOvB0fsUjBz6it5w0nYXfoZ++Qs
NVxuwQmvvNyKaGM514RZyddFHGat1ZODC4CVDuDJMZ8bgP3Wc5i5PbKQu/+Y5s4Ep0YDMqNEGvS/
TAmBvi/aKB8R1uH/kUyOvbGXpaQVLgGoTY3j+BIZFsclIpiBQ6ne6VQ8Chgio0WPp7qAcKvOvUhL
/yZwOQXYNAIFg/kcKMcMzLsYQ7CmrKQLIA6vdHHIOJgLJg+PegXmqlNOpra6LDKptZUADKwb/lAL
CGkARs9bGFQgxcyE9oAJvNCHFCwdfVD5fk/aEqSYX+VRrOySmibWtR3nF+omKER66/ccgyFtUxMa
vKQWMM0jrQ3sWDmjz3H6xnKHsztcGHN6gGlyLfIdh/lYsmQOz7LVCEjyXeI4qSZ+CkBdAwwSf3Tg
qZcgCOKA3LulAAbv/4gUoGamiAmmY4gbtnK2S3O3XHf87G13Qk2FmObgbG0UM/y+3aP5SR+qSMNv
ZZb0JQm3mD3wTtL6xF6EmsyucDXJ7eQZlM1SYtwbvywaFliJDVa8Z3OcwsYQHE9ZIq09qY2yAyy7
WjiDK2Frt64hp6wc1usLD992HIR/B7Dd7ZmixaiJ517A3mBlI0kEduniX9YgpKprW+t8H2WRalzU
jHE78qX7NZM4qIYRSkrVCGtk55S3LOC7MwXQowO5Rx15NP+hoB9FIO1voOXt5qzUbibZjO9Yy7UB
vwVGqULNR5pBotIiZGWi/SMUGQ6+n8Svbwz8a0Uav/qmMU+Ki1QxBAh7cyeTCUuB0dHNjx3srTCL
b0likBf5JtWLnGzLdm25kEnOXClnTomg1KhitFEmeumaQiN7wcYgq19LfuUXGQj6C7EOb0+H1TMh
R5DIoP2tLO1GZU1q2XN8SomDFagWw9Naixy9AAnSTXWip++EWguXu5oCf9xHyVH1bG3taLSGBAQd
IclY0O/+gebj7hjUdVVN5UBBWzmBlAG27pMLRjZg4x0+eVv+lyqJg+1CVVtrVJDomTq+lH91eaOT
lvSEDs2epY9oK3QnDvw7nVOVy2kqeMShSlaLChgW6OdWtU3XXu/ge4kjmJ+nrgT8W1GopoR5/Aea
8xHxwUYcJMlnseDv5YSaSJAQMpirZ45fy3s1NHTqmmNZWBE8Scai3ANEl15gTCWXuNxA7Q4iNj5o
1dAJNL1ZRJi9AKoWBqbmNg2Bgjfsljbs//r4jY8Fg2rvk3ncNDMleQMCuzS/LpI6BoD5xuga3DvW
kImTbBjT/ZUFY7jY7IE2D9tLbSGQMO9g0oPF0ynd41Ujrhkne0mcZSghMdueHgX3OdlO2uVS1Fit
dgZcAe4D2Nb7TL9YDqfX8Pe+VvuY1NkQzTGzDtdXuWUPa+c2pGb/QezBqlW8enbgDWxC/rR4eXKB
VqAJCyih02aXCJqTdlBxOQZXHdyGpDh5aQ+I8dvDFzjZfiybI9RDHHgp7WJc3PMq4KLK0icQCs4t
eWPm3ldGADA8GGvpmHM2GtU5sTnZ4mldr0Rhk/BbZL7Mg54jd9F/45AhgzRj3cMWkhkzldrdW4cI
0hOIfOdt6W7joIEo3wNFkoc9NZHNT5bDlNuYMsCBC2UQ3GcUYdAj4sF/6bRoOFxxLUwSyLhUiDr3
vydMVKWhLVC4OQl6FCyd93CnBgZrs9m9lNiprT9SeUE8kHql+rnJ+/v1HO/h6NgEC3wvfGS8kzxF
9VD9MKQtHB4EEdDoomSSCRx/7OZGOfeOh9nQVOo5YzST+SCdEYAwxuSUGrd9hOSMFkYYzytUz1Ah
9ODK6nvR/uYBTAnaqxQKC7uJGB43nLoRsTT31XEDTFB0JPJSwTFar6BTgfEOID0IfzFarIWXli9Z
YL0bpiWUJPNQryuQmkT8iH3clODY4E3Ezv8qBhf0mtlMmG/kMSO/6FMCD77NQxLiKoLo9Bmpscjt
8UrznERIRh7oGRWFhL9qRt4hhF0ehzjxxJzKcI8VFFskjMjlrOINPa7p8CBErnaJyfE3JR90x1TE
3PagMJKvyv72hoblYQWeP+6RazuRXLwNr1mI9QDyIJ8btQ5E3xZvGYjMwkMdtW4kKYQQ44mABD7W
DCdgnz5P+D2QJhSfMqZBMz/MFIadI2pUOFyXf8fvkOMzp+0p3WZO1d4e9iXJmBXTjP45WvqhDzLQ
DX7brQ3Df2x2y5efcRQrVcpIN84beELjhq9PQsxOP1I5RglRnFCJFjB+j8YatafpBGGuqdOusN/a
jZI4cx5ggNoah5dGuUzmuqIQPUzD7ANhz/3+1Rmq9Ez63Sanxs5Qu3J3FdcsrD+39PlGL/mW5ONy
824tx5MOtwdI/arV3vJGM2I1zUIeyWfBNreZS422CriqXQ6XnRkLUon8OE/VvtSF4PY2ASMRlW3D
T1maVpVShn6Z/teKTAA/woCWmUZWgIJR4OaiMJ8sGiecd0G/MR/KpMBjqQP3XDHgzC9MWZRmAKNL
xEmQXPQlU7i3OqyjhtRtqXk8H9+CDy2FEIYbdebO95VMEQt0yAO+1y6xvbMZmdHiMvwNkyyTuu0j
7vf5wCiXMOryqfjBtUY2vUx8ops/QpnzL+CFGCqtf1vCaT4JPscU8mbWhnjEuLIkHXI1r43/FYsw
ux1H3wohkXSsy6g1v+GiutFwPs8dO585UYuJ7e79ZJpClljejWTit1UF8vricXzqm2SrznCEJbny
XQj+83TL1SlGddat3MmunsUw6g3D059sM2b0pTyVuOH0Vv46iNdOtoNyoOm6hwA6oFka/XTpHz2d
4jfh987LXky6TC6hIfpNfUPAOgCZvCw4wqMKWj070eIOGWDo27T3reFALwO5H+w4CYIb7IV42JtX
GRGyFYw51xGlHhZS7QU8GFtbraGQdYXQPF10LJIvHnVuPITjHwVKv6j+AApR7kb0eYsw1q7HpXqo
i+lsqIyCOhGCNhV96gyh3YNoK/eR7YMDYx4uLbFScAlbWPkWFVoYaeLo2DlqKektxpJyOxb4ziCf
dRBnoplAHvvspzgHVoSE7FGBCHQ0HwVZLiaQW5EqzrX9YFUD5ZaZxEx5A15i2GV1f+3XLEdXFRe7
jSxAuhMgWReD1NtKVBpxccWhG2KglbCcPISfG+2SQLbg3YjWO09SX4S+4JVgll+5toRkLoye2tUd
LXGIl3GA1RlYS+0rIZ99IHK4+wkOUCaXV+/v2+oXXhlTI9fRzTWiWfRxAUtZjm+RtVaXuw75XPSc
gcOy6Xh+7w8mmAETJKBkx1X47zOajMsGvNSs9UJHEkp48demgM104dSvEQ+RgQF+TDKiCTrZxpum
scLOoUa9TFqeSuXqPNHC0hkklREpmLg+Znt6rJZghk+RJobSgWMKsGmQ0njUtu9hUJp3kcf08bz5
WBxaC5+lToCZ8xPGJOIGWYdVKnMvtNGU9gcYQ4K4U976eGekoNmTfWdvl4UGsw06SDn+wPOrXkjw
tdoR6ARXuhO6RH6ueZdDhJv5oLHYhb4SFCDKNUH3BZdqNmRUMhMFEaLru1G+lWV1eFmfYDuYHPl5
Xn1qmhEcEFQRZpmvrJbi5hoWmqLmzkAfbZ+bs/Kb/ZTSKMFn5Shtck89psbygm6YexuAf/u2TVNZ
hFxnV4BJVuXXGCGCeOT6W8twatTFxr/r9GZmSIW6JA7UPg/360vNzo9i10aVbTInzEkJIdm64eRY
rPSddnCwhmXki8QbXfkwUj1fDK+uIVCFpUJKBd3sn4eFkIa6PfUt3uqKiqygx0GHHkdGXVSD+cFA
vvf2fZzpiRr7X5tP5FbVkiKIUyQoaGxiGEnfCHhde93wZ+3RD+a9qmpjeKS55EdKpMj+UJHoGlAW
9Z8HAH2C6pZfJeytMMNyEpKXDtsPjhrjc4MpzvMbhgZTSQQyBOW635D5n13NMa6Wu/eYgbJxJV7N
9ApsB1XUaJ6Au/qlJKvmFNhBzb8xNKfDyKbab/yK73dOsmOt9dMKhUaBQGWd53zUufcK7tNH7tQt
paJbVpcEVxEIPJFrafBihhH0qx+YE634IH/3nvjeLTOX9/96Ix/CEJAJpnYJKnQ24koWyN+tGrS8
PTMlAyFywfwuoQZUNAO1XW4PYxbEOzhKZcVgQp0sBvC0ghW14SVjk6P7qbRLaOTnxyLjn9rwrEd6
RzKwZOUPsVesgXD8OYKtzZK/+LEcFj+8XsSvnRRaT2dtXJC5abGKlqKOpfqslR31ghUPMUAAdS6F
hEOBvSZgUox9ZwPqhnUMbK+QvyQENSBfDuGquc40rghWA8g9wLMz3q62OMD8X5L28TFBVKH82/nw
k/nVyPHKdAifCDjuVICnEVFAsO1UwUdaLpAIMrN9sq6RjDrT8ci+nRReEpVP4uH5UUzWV5RA+8qr
0Dj6zJ3V2sq23h8XMuU6Ww0qTq3iXYvFS1kHqFwpWINDHQlNZ5IMbgw02M2ugAKDJo7C0rWkv3Rp
AToARcv8oS3MMBW51dSZlMmUo6Jkx3R656oDRX8lH5jjIeSSppK8Ff+ZjSf+W2fx0/Bbycck4a36
GICjD5G0gDBZcEWFMr7ffycIWJ2IbaILHzw4j3R/BJh1CwpwbPIPupp0dxPHo/j1uG46IEAwZp/v
hUzaDha2L8D+u4UPsSekyjbOwjsgy8ukLyyg4EbpY+3JNC33T8D5w4ftQ3PgGv1I7S2CCiFUB0xs
f5i0LoAccvDLMFHpxLL+znb3unucLEKf+yVf8NPmqUKX6CceAF8OBfUoi+LpyNUIEVh/ddVuhzkH
xi1HIp3mQPs/7VOlpTzDYE05sw/0ob39oNzpG1HG3w4qnQZw5yJPnohoxx3TsR/utd5V03MmB9w2
IcSIMm3RoIzkyaQ3+r+GP6QqowjwtNSELiPG6VvBlHk7Y5OvwIMsghwJq1GU85QABssm8cwRjbbM
My2zaobBGQrDlGpftoZkn0jObObtvHnDXoUGsr1nTsc+RMIDRASgvUUKfe83VT0OfuPbVmijZJl4
jrjU8nj9oT/cIz12MkEV6GXEewLIiMb1iRBjR289S8IGkdUX/8W+HmZ9ul6Mf96HYXt9V703Ek7P
poJ9d+H7QkBdwkpaKIuUQufDFz+36jXwHJ8k8eQB/CntKmFSXLBhwPQhSIZUEI5w33h5MjNx+slk
DBEFh1NaVU6MuIR1qdSiRErIoPtiwgJjtIQX1ZGdPSESl/2yJjAvn+Q2z2W3jnpgChN5Q35hxQo1
GDWAhWMXwUxf0sKs69x0LcSmeTP2RxNHvnOEJlji+65KUH4IpB2lvo69JpuosBmTFe2+smgWLP0Z
nkL2zAd7BTwcO0JAHK2+4snGrNtwO/Q3DdfsNptUbziCiCVf+f7WlNlfqGjsOpY9twdk1i10ZUml
vYMyuhwkveASYvfclTuyfpMO/a0+LETfD2cR0vjcdE8V99zTDxWfgo7/trVPO9V+BSj3a99yHSJ3
f6lNoqSMNqnMzLfp2pKcgFTkPbHH2zyixim6P02Vbk9uI1mCsoJS14MryM5DF+c6yiOhcWLlg83z
INI3LNB4Uk/aEVQ2Vtz229bFqsUdjW2F4teoHO6yIpd85gWBgRK1zwXmJnVKVDF5XyefYwHJt1qW
1OhVqVIF1k8NTYhCoA+QHpQDCXRBLISaZwdOb/YPoDwJ8L3KFRDZyEufpxrTTrrV7LNsKfxwor9y
msFDHK0EILfBettZMBdbglOuA4Uu1h/iq9/2vaBPJABxxPZsXn/9DibQv9ue1U3JTB9lgVcWIW18
CkERm20of1B9syAdqIS1OLKn7pf/6/Z54/mxDQMcUMZMqjOYhORZQZ0nGfCDisWrazjGWUUG73Dm
T9l5caNl9m5dNe8YIt5YqllUHiNs6lAMm1GObcPtT7BYbD7s2QuMTGdS9axcgU2kbYHSkXoY6KZt
/F5sCxoI+fMW7SJUAAbFWwdda/ipc91oCStSO3UjjOTxN0nCJt3iYqxZ74stC/sZVDXhudxuq2rL
0B8GFAnRhhlDqMpsfWWfHxzc/jdE2aD4OhAazaU7+7RH8hjk1Od5Pw98I4Rbcop//XuuRC85Mp32
rEDRbnQkE9aze2JGQRi6ke3Rrt3CSUjvvPlyI1BrOE41DxjKF6rYUzTYEw5r9CrKUJ9HLwqx/hXj
JBF7IORO5iRtW4BiV4JwzgDKjig8prc38yjfPgkwT/xeucnprZNJiKE+EQ+/kfRHpFfgf7hO8am7
DERgdYB52I/0WLJOLDYztAkdP3I34+5FVnX00QcFJQqNHq1MtmBFi8xL7n9IDa+czGGZ074QfVlP
TzbnPADM4qgGiPhQYL8zVh74+ywfpITOY9Ydv/f3x0avMkQn1o/+V0q7X//D8bANg+5Fpb2brnmz
9fkGDYmbSTjfJZ6cj6juby12DEnHJOXn8b+nB7ys/gv9lt+pWT1w7f1ioej5E+l/hgNdamBKbflN
ul6tZcVNHJz8FTS/A8KXCqOljZTFJtSuBq5KZuIPx5N0LkSt+LR2MBBe3qwjEYQwN546Yf3S67X4
X6FbgSiWJYfrQ/l2SYQEs1KlNqthHgDOz8S1liERuGClhmukTldu3boTJwephTsS5r0tNhQ8zuta
sYU6XEmmPav6zYpzBrkfyO+dZDKR8raVw/ruilGLJJgkyD5qyj5jMmwyaMcvfwUCF+kTH9AFPnl9
JZ6fGRLf16Dcsnwy1+PE6jzpDo47E1Q1SIFxdad9KhOAF5wI1tp6AiVpqQ8nD0t7YumrR7F6EGuE
7wIZqGXBAfzAcCg6KDwSXjJ4AlATJcbwb6W88iIGzckAFxcMR/wOgHHUF3N3684oe4FDmLuhwr97
BYlc31M50mJOFC2GuP8zoa53lNgHR6bSqAB44uVE3I6189vzBjXsJaE2MQMdN0C0kC3aQQ7UD6Gm
JjJp7C9Dd5gCeqdolTKPmu/sESXA55cqY0mDqzJwEuchHAqkJCdHdPRVxWFSMazqWJl08NKKCHdS
Qy7DWQNa3o9wTXYItVU65TL/F3S3txUKP0aYs4mIZMABw0uCUXhR2d+d5bUjcMKcokaQhcfFiGdF
oYSAIakO6drnvz390whbztoOmEHmkWGrlYyOPSxNdgrAbZqrjrJYnkMpAu2Lf6qWgHs1J8lH1MOz
L7atchaeaa5/BYDmwBRfzin7r9/fA7o4OjdVnDw20jkwN7DuTjmUQhY+usjRk/zFlF7NZQtsSFuU
p8aDIiH0EW11mQTQ7IScPCBzbvW6xe7X2cF84bXuuW9biD9m6OP0FhmvdI/OZ+AFRtFlsO8mLe52
5eYFXhk/AFNZZQzrxXnVJ+2w4OYXQj4b7BNUhNRw5lXyq7RSqJs7iwRlXpT1O/FEiwQCbjx+6QZC
WDtTk4FC8jFVKCXJ/YBCHJVj1USBWGgP2BMfmu4Jf5cYXTX0AEXauxTmUIm0rmDhpVxqB+qpoeaz
tndKw/eZa3KkYpm4OFkRhu8PZka+FudWr1gHKMGSUuepv0Rmf5xjcmUU6UGWwMpYjK5m6bjJqXGv
pocbnvhCspYB6WBztrKpnykLZPQW4dxtFGa4KSVAHUBtI6fynMwJeSdFe4giYMBb2QlYcIWhzoC0
JFd85/K32/Z7/Su6ltmPvByfKpt2/PLvIk+lWWx5D93Tghxx2Qks43rc4C66uldKjlnesg8lmgkK
GCAKwlMEikjuxYmVekPALOtn1b/PGuQ4BCx3UIdvgjQiEaFjhMJP34MwrUd6vBi/kNHu6pr5xMAS
j9dc0Sn9Xp+e8mx2yEZLldoRsXuveVOaZ0QqYVAQyO+GnRw+W0Iu1pRdPxE+aNrY53m0aBYhhlLr
zlwfrucMqUTc4lSu1Vjl2cc3HMF9njdREz6I2bAH8a0TRXFrTo73MB9zzd8xlnEM6bVfebziuFPa
JhkbmB35EeBcGTvQuNrqVEmp5GPAe1Ih65sf0O55pjCPJITU9q7gicSCdtknzciwFmZ4CgUFZvxS
mDUZK9L+6R4gv6/b4k2TafQBzxohEG1SF2g8MVNac2oXFiqeMwV1Jmrh3mWHMTFEAJdrrY8mlq0g
tBm2tMBL8d1g4bDf20NfRAUR5RxQSoK4brPjvYzdyKf0dfLv6Nr6x7vTQHKITqnzEDJsrRsfWDtb
VRtJkg7+yGrqkwBEP7ELe31oJaDONG4hL/YLciW4lJdscI7NQIJaKaj5tpl7/2c2ua+s6OjM6XJn
tjRuxterbjVGkQfmrqC8kNsZeVVb2F3TuzyfczlQ/Mx7SzJNvCia/u6b2+zvg21ckCLg/Dqi8Dyg
jq8fYzc6XOBHnbcVTG2yiQclxFsOQDyXnjkX/bWNHhr9i0hZQufZdoV23Mg7+4plG1TDvOZwj9YJ
pw1yUZt13KhyrcS0JTMPLiFTmndZvJhxy65k1WT4ScBSMBB0jCH4TsN9Q2l29aEBXL3WGsyvIUmY
5I9qt7zJvK+JnD+RFxTxYgXBX67CfSiNpBKnyKZ2RCK7ItshuQn0bM7erxMLDNhWbWEHE/G2IkMO
49w7Nq9OXftwiakhA0fPWsfloXG6bVhwrvWQ4wIE1ypCN/5gkFfb5dDtHuAxH/ou4eg3VXUPGN9A
SncIYxh8LoGqjgXv6aqqDBa37mJjrHuUPh+7LxteKoil4J2PJB7c9dJYo4uqe7SB8neMu+uoRn1o
PeLFA7gWjNs5Cv5llI1IkA1cv6ZHSXCLxFfpidu06flP9NUYkHFY4P6gdRnMkFMpjghbzcuk+dYq
BDhSx69RF07nCZGRpkntFsKtCj+5XbUteD2GZpb90s079OOLb107PV/eIBmoTkug+5zOiuytN2xT
sCfzrY+ByrMGg16IbPIChmqiGqyLD3Clk6eKZiI4jnRGANaRYPPutOSRcAL+UvmpTDyEz3XAO5T2
sqjdza1IGkTsuPHmt2qJh2DI1aLqw9HmZmxIcSFBz5usu9u1JE2Xg4QAGI9xusMKUM8WxdYC9EQi
4bx4Uv7ZHQQ5ktfpMb3MZtndeQcL4qmAVAidLs3g2NoItiq86h8d7bOXnLxLFAIOtTMRvfzBR/2Z
azuCgevJirmnKl/9SrQQyD9zY9lawkAK37m4QGeX32cdt/psm1hftosuclCWr8sR5O3loI1ONnEK
cl/lOAbETd40mkgXfcudelYwhRNnrv7h7WKjk7TzXlCbGaQcr67JnOZduRxdrKNL44jLckddN37f
M0lYeASYr+4hpG/G9jCi6hqV2Kmp59MYwEv/ZJoRlPURey1+3RUtRHESsCN7nMgAhnbJgqu3axKY
XmvMJzRBLuH96Eaqmz69TOiM42Z/1BE/d++TeLrQlh4MmY6w9kwL6P4gjtb1EAiXGDc8hsvzhaBD
zAjSrYNldJH8iTUlazLr/ogCNG+IzDl3cmrnqNbe1Id4JprMBEwpopwuoNEQkgrhGFUL93J6qQLr
NsQCipJ8n5P9TE/TeinPivXE4Arzbw1SIDLnI3mftZXTtQkVPEnp50kuQo9vn59cve7QqIv6L+XH
baTKMtHoPIxUeZ9zjMr08Po6HqQayYxaMf4rKgQ0HpjprjbYsoPBgSrpurSNjJB5LJQLnfj7rY23
QsDEj20/LswjzQVV9dLQuI18GOcFLVVERAmsYp3/GZC7SCgNsg8TXuDYV15GSdR2mgb8+oESjBev
mfq+u+ag51I4iM6huyo5hNCo0iwC8Iz0JbSSBMg4gqe7JOqdeTmW4ekd7KS7FB4BF7wYUn9kF0RT
MwcSTwyU5lXsfE8Ry9oaNvOxrxyPaOId8L2ZuaR/vfD179+dY/oWPdIG4LaVAYXvfY5cTSMZNqPu
YmS7rnDdzCfQpSjNG9b0Ba+T/ThfVdbvDM6hQ3whpKdz7WplTkjql5gva4BU3Hq8v5akgQJuglZB
21qf5/ZzjaDs/wLEN9i9cLHmfA5w7I69xqSa8qRxevWo807/ZQineD/yt3KA0Qs3ng0TyFi/MpXC
KumBW77//iifl20GcZyElL2DaldDYv4HSagT59vleDRlY8ouWHvG79Cz1YiRRCc8rvlF07IEdr6B
wp9L1VBZzeGyYBtKfipfDEx4WPJ806VJNz0pyFr/5hbM47X8omsIZp09I6zCvu0Cld15n67RDbdX
u7GKclbSzyA41M3DRMkdOd4ZH+RMenEnxIvhr9Y/pEd7CXcFXkfgro98TD3EJVd2YrScquZ5jSJh
rWQ6i00lRELL+MMnk/Tt49f6nhGei7R4tECS6Ygmrs1fsHVV6USNt7RoFYhcWcU6TzsbGaaT/WK0
/j3x/ypCv2EmyZ8ir7AWQqWBiKUNCxzgrQdnpCthbDeaHB+8I5/mR6zsTk5PKVz21s9o/CoAEOBa
yXbKFmViEoykTojn0ty65t6uiz/VbkHF/g1dcO7i8XDoa4O7lTDoiHeT80etXH1cNNz0koxniNCe
4e7lkJOLC7DvGn2vEOy0oYdRxLKb3uqdyDd6VI6zCcGWZ/9jlHpy/1nek0eV++jfdzTlI9CGUtSN
JDF0ZdgbbbC8ABmpMDONqvF+DVW3gFpVGSpc3UJv80ciFcmntCl16Jt00dEtqcHpcaLIEs5hDKPQ
CBPUWbO8oFCKwNnMuwQRuZ5DPNQ2iJhQpzXhCCArZcWbOQEpH1yMQ0cgMNPDYTqYGnDIDhnk9hsH
xKgg0AWc6isF9fv6WJHop2xsjk48nBPknUoEIj/MDHxXNHmmOdtISgugUB28dvTYBDOkTkx47Mhp
uTfpEX+mTQb0Jaadj6tSbhDBHsmt++6opDzvrzoUDhM719VoUPYbfGyLmznGarAnIvc+i53v17ZE
gZ36SEQIi3cs5lLsKuFLD2W2u2dE+jMg5G6noAG1KIEpIQ/OkrVngQbl7kObLHiA7G352dlWyJqg
nvgc197BIhSMJUZb/o3EFclLpwnTwZ7lAEF41i5z7Gpo9c7Hylm05OzFI8Mq8cod2klqZ//Nseri
0WoLUE/TrUQIEXST7V6NEXpk524+QH8QymHl4PKI9+3E2ToiNS2UmPlyswYI1LFd0WZo8tMLVUXN
kqD+iIug2RMS2bhEmbxBz9bYEUedlrR0tM2N4RzyM5zsozHCT9AcVF4R6Qg92D377kiD7qcGOawV
R9DLiNCpZMCcW+sz/AYnl3jFgcKhjFvZgWoJa5g2E3ouDiiT9pMjeXHpQQe3+sTB9diHPcyq0DOZ
HSkSNn3hTU5wIJAc+N3Gs9kwieKjJFOUMx37pDcvG48OSNJUtn2yq0tgiytYT/TxUU/c1rhBEOn1
3dD03ye4cSnSWgjV91UApF/SzQaZdeu7Q+l8Et6yJ35RaNYZ2Pln3lzkhG3spiWcOTWaFtkOeLl9
JQ68KxNYICOreIYwTBy8akj2T8MRHctc2wzSmsNMm6AhV1Vi6QdVEEUpenLAuuxLlKm0hsoeGdNP
ctaRSuVS8X3FYa0LzPrAnSpjt5xCwoaNt2zatZp3lCiXZGo3YpVHFQ1AJAJVK4bGcJh05BPEPxYR
vvcBjMu/zEDm0ahTYX74exDwYyYMX/30l9PRsZqitPCDOjqLGFZcZ542MJLNAsv96Z3j4hNqBiAY
WHvRj/cxuMNgP174oU3ybviXZtdxHx2TNHo6Z1FkjdxFPJzuvarvt/zKThhko7OMReB7VAM0QFPe
wGlfQztqxUgbUC1Dp19Qdgn9UxQswI0MHYU5o7UVSNKAr9YU7iqtW/E37xW6/hR9TFTB3sZBrW1U
RR4DKx2RZdZ6UuCCiRIdr0bbeeV5vxBw9wvsp5yJRvnrijYqPYAWcK1gYioz8u1JwkkudDBNrA7J
OGYpzBtsOL5G3VXLdTFOrzfgshsWLxxrTjNNGlmm6rWRb9AWu/Cfw/51eYHyUZjjV583R9htewLz
Gq30JeCgFVCLYIlwrTb9vqDefq4yy2Vm3O/J/XsznXWem+4uRIukfqu/fHJKPW3ECAL+zWjEupBw
KNH4VcjJ4GWIdw0cUYGDNX2q3JX3IOClJOOJ3TGVqCmzQuYXqg/xvLGl2G0BKxx+E3UsqjySJyrp
VG1vEQkizfqCmEcMlCvho1PaQkCiL2VkkTdWdW9KEtHZWjQPdSqRyMVn/ITn9RG4SLVDU4HGrhij
IwDNmY0Df5M8r6Xe23ytsuEsvRpveZDWd2S0YKxpOWaifbPPLp0NUNApwc8ZZefJiwMQBYP7IVE0
XIf9iEBwiAYYuLHtyPKc5HCguu3URHrI1cnNKD1YSIjG7lnAw7ggJyOB+xSp4qpy5O7AYDTDE8uS
hgrqDa5a7c0DPOGUP55ZrxtlC0fisan3DAhlVraGgkKTpKuyUCteAxArlKnUCaOMotoE75ad95CI
2Xijs8EgUYESuQ0lN7r40cLK7npVmnEzdRJuMn/cveGG7uqmJnlCxpqzxngOWkf37/2paoztWno4
b8Um59mcKnZ3fjmmnlpscOnkHIhVGPNQ9WgWE1KKXj37/tWRjlYuzKsylyr8TAO4LbEgnovHo8s8
tdEeNAatUZKjn2CEC0HATQhu2vjpZANMrwhgJFeB1JYiFfj3kF9V8AdP8FzMR6S3AJ+AUp1BswRw
gRGMM3yB1Xq82D88tsBVEyfBZk6d0HVXrx6tioW5DeQF4pQ/3r+5W/m1Vby5wyZ3q+8Md+W1ejLU
skfBjBMRKI+WlSjY5ObHJrkQu4G0SBUio9Ye88yj/WyPwYugWJJDUUlgtZdcgJihrS/66sOMrP9m
E19qBsEcyg5cTef2dmq//lbtsIKEcj2c8cVVqRWBe4H3xwoHXEDxYr+JxBC2+kEO9DgYa9yaS/7/
wEJsGDfhuDysVz0l18afxJhfwIhxFfI/abIo2BlPWePrUYSBidzaW6rOsGAfYdWlAkIAu2Qh8vGn
vQq50GVUQPJUGdx7Wb3m/bJtL2yZ8m37G5iOqGVE03ZGYB1TRu40orYryiaxONUagZfrvCxSBN8g
tNaw1a1V7HLLnW4xJMXXsoGSQlNuITQL1NZVI+D2WiJsWujN24Ncbhbiov6cIkVv341WyEcqrp4p
jCWsfM0X4iTSwOpEsKaRNBrESzzot6ALreJp9IsCfsQMCAlz6aP3yvcG2F7/A5iaMZQ1R3rxw/sL
sEGQWZhYeJCFEslCDp2KosQqNYWhykmu91mNbUfNEFM5aGTX6VQ0Xtp8XDtjyzWdGaImu6bqKoJZ
Wh6927OyDrjPn4VnDu6qQB9RFrf35XWj6mhdn1bICEplMTSdhIM6nuTVg+RENQxp9HbRwqb2DNXi
KYLCNllyC8jfiksj2qWFFu2AtFqX9yrJpwpiP+q1U2n3vhH4fxt/oTVZ1M7FEYGkJToV6s+8id92
FdKjSTx/pcNRC1gPVH8zMp7JVyqL/EIPW4KPpv2JbfjaP6eg/2AnlrWK8hIWEOFxrZ9YgtDnUh5u
dzsLd9iYhCMfPxDCNnDJUUFGfszVEFpQjj63ePsoKKngCQCWvcvRZS2LG/A1WWl05E99Crli8JQw
/1sAr5RNeK7tim9WL0XuZbeYoeu3WVhHNqwhQeYpjr0dYjZWyv7eQA7Xbk/lJMtJIPEtZGEIhZmC
8dhpLLV3oltHtm5RJtTz7yeQ23eZxo0jflr4WfFbJUif6mh3lf9iRhmroIFXk5EGKiN4NqHxmQmE
6q9HgZFspyLTD7uNb8glDnqbLWuoYNig2zu26b2lC9iE/VGQrI8MPB+wSw1HFaY5mJMXaBYKxFeK
zra0w9nZff7E+J3jLdFqSWccFYGapJYBvRwxRBIwGw93tVT2stzWM9ZSyDUtLTenoS+EXMTqnVtS
0n1rCM52sTnLmB/V9x3emrvAIGMwQchLIyKIkUkfQef39YYPNnkmjlhg7sUH+7tyurpJyNEEC2uC
qPf/CkUDNkYGnu4lx4iqNokLzI5rF99Mse9pGaD1zSpPVPdpBOC2+8VBOwlSxRhahRLW2w6MxiHv
YgMiUkKgyJV9Mb56HgcQ6OKt6O7wYMjGTHoZUt7sfU0c3ZUlpMYuZJOeAacEajt8n86qUXJesxzK
vbiKCa41uk+ssCnghK4U/G5SDfC1kZEWdDPkGnCwsEFbiLuhU5OWSzkgag9kFxdTjYk+aJxoGGLy
oJGDwsSKIgIY+p8YkjbLrJU4oy+J4X6J3YkT2zz2ZTbcfKxb5KfsaAEC1LeqcLkT8xI2uEzW571t
GojTSTTNo9c6qTes/Aqo94qERzgbpQC3ODSx2Z9yokebrZfp4AJOYyJKIRjG7F5AJpNGREhFWEHy
PL4a6tLKfefEvqyNWOEIZx0vxAYLCn3EDTcMk6I40v9+ON97kUNSrYSCE+jr42GraBmE8fNddXhh
ZwCTdAl3jeIqHhaFeggjDf7b/CBmSAAW6qPT6A4uoklTnfQlvyFCgjlNUjWf6o+F7GMxnPp1EUmE
InRDhLfJIpuiHCpu80SLco+5pT3gFtVDK+s+pq9+6KRQafnt2Wt5alKvmOIX85o0ZvVafvSMN2GA
o914tcTUJR0XCFFdkp8kvjt2IdpDU7/L1QUpHjl52OJNSHJ55gV5VA4L9sgObA886AlyL/FX8zp4
Ghx8d1vdYSThfOdLZRzqc0E9A814eC/EYmnb2U0ZCGdCXmwAuoc9cnWdXoMJ+j8l3H1pK8rVazDd
VT1OTRd74OmPXJroIb+rYZB141zFMUdQA1c7+ftO5akvcCEGIHlEoCIEIHeGhGhu430v15+a6bGn
UWrvhXuBSlCgYfGXszRiOwB+HbtfdUDSoxKBEYZK0NTSOFbzeECYbWG0ykavgI6q/wwlbE548uPF
uP7VkkH63ht39Ke8aK/ZqQLel9JJywPc7OLWi1lf0BxVBL/mEd+42KrfEFZrcsvkXnr+1Xm6ti/Y
RXBm3+O1dZBJc8yblZ06E5j7AuxJhlOMgUTyCiSO25Tme6HgANFQXIRKnOnEAcGU5LNn85TjUYcg
CX8Z7/TfTUE9xu9DJRmDic9B4OhF1ab1YL5eAbq27PP+kl863ZCdGCw7OJfwwIHjqFNjlU4LMfNk
nveFFcf3lhFFbvcPSIt6Wy2iHCrtKFZL5d8j7UDX3g510iFdikoNHKfOUh8w8A9TweT1KOMyL7aR
rAGqIGcXa7+b9uuE100mmVrNQJBkGex8HrYOYBDqbdLFWQXOkrwSfG/N0Z1lSYg6+7DwE4Ml86SW
UexVoUhLHNNPtUXV6zQswrkX5syPltd0yD2O/guj3CBEmFWhSLtrbBEozQEVh02uIRjIXY5pWxgY
zjzhZF9S+hsQiVFXlL+zSup2qhmD//ZmQfOVyiDKaCqDZ7g9k5ttbV9oESfDXL1rL+9wzJZmfWG5
nxm9RlJ89AVZJCk9xXtpZBvafWooZbYKn19lybjs4tBWHfvywsguWJ+K/gGzpTcTsImeaYAe7VFc
URA0ZkPgj3QkRLXViSIiEOuE6EUEZHyHrwPg9G++Xkd6PNi6li2M11a/gkx90ZbAc5ckhfSTetar
87z5anbI4aEsx1zOL6bzT0apLqSQY4l6gp0GzYOqLOWPlHGOcgdxdlpl0aooxWbWRtSS6/TtigLa
elz0JJkLg+qNh5qTRUGwZp/07ldaSPSgECDsIWd2a2MZdaTTU93iafua1zzq7Z7zsxkFFT8n11be
tPxLznm7KcyCJ6Lc1QXGcXiRKpjFy/nVyRL9r7wsj/wLKnjfVFfAnFDqSeVkIu5JOtnQywvBM6lb
NM3Eu25yEvAOA/61TfEePLkACwtH2gQkrqLsTxmRHYINP0411Xva4Te7akR2yY4MRdNB4eXHdQYz
EWvCFb8QBolDwkl2URCSHJogIbCI7emNCMZfTn8uyuh4bmC39CgK92PHUyVmrLQrtjYosI0ZUGmA
BSHzk52BUZJIcwlvCl6Fk4EO5x+R0Odg0EqPkljK/IE7mxyuoVPGqTZ/3jQpUpi3h3kmGL1YgBpy
q5N/Y+n0ADkFNENQuIuZq6cL7eXExWYy/hd4d42UBTXkw5p501CMqmyG+7D+4SG0GZv5+xLm2cTu
M9OiEBME+tiF+ZwhbsCLWT/EDRmw91+TDZggC1GE6PAKAsCwNA9nmRsm/KWf9o3JGEys8eBonPvm
rYjmUaEorn4LfjuJe8/BeJWEgkYiaD6VJvwKeAcokvBzV5OZPc0JsYaHFJKtyyFXvg7q652qEC5L
CzDzk0YEAA6OQ9koQ1etWJmK4H90Kf3uJLpc/+QAC17jON/czKY8NXQ+pwXtV9HffX2nZIr9LcNo
aCZ8PcwuBnVVMSKrQoBAHqUz/+zNNyajDgZQxBg+XqHuMTRn9bKZ2eGxENXQWzwbDWiwMX48vejq
grnfyYWzwdDMrIyBuVXh91MPGmdiJwMYqxE4SnHGTvtT9x7T1kuvnb7AVC9nvJOU9RVm2zxIKPOb
DagUywpwOoD1vPMB1uTgJ0EbjLlFneSkjk9jKXuXRNM/OGeTXYK2V58n9qirKwsblUxdys1JLm+q
wgMWAUWeXc/wVlbYsMFCk6t/dKMZiXTr6D4jbhNFY+xKCDOroCEhR+ErMTW9qcalMm2FwmfTkAmy
plrN1lfEoGQX8whmnkUJqjYlETnsF9nxegoq0ogdb+Is1+PsijqVlJDKahKibGKvK8zy6/sQfXWL
j9QfEHqo1gk/KTjfxFCCD/QM21kVLfLKQA2CO/8sVXxmk3obBGa00N3YDcyE+U3gMDQQp6nmR9Io
vqqLUDj2DzzGmQAPz8Sq+0emxpoDflEgeZyVfke4K6Bkhp063cWqAMIQavKN89W7bWGq6zbXzKFS
MYiQPt1GDNe+q1Lc13eGBaY1PBRbx7TEvLK7KuYe0nWoKzr5agXojtRI9akLIsrxXjILGvecLBiJ
onfHBivDQ9/uwS1dgXJIBzlzzXfkjJcZJ+SIJtBhi/PN7rCmkNeJY94eLiyzaOWkaymrs4K6r4mu
btDgtxsXAk+BzisZ899QtayfKL4ivEw/w+WgxS2nWVysfO4hAhJFsLqOTh3+b59dpUc9Ii3Aket6
ggf/gwMnAzJEfQ9tfrTIWoQHm43NfCcPa/4z/RrXCBjn9jhDL8xXUGxyflD6WUAdPE33MOHSp8PF
SC/m6wqjIudVNBpfkX+jO4BvesaCBqBiQmAnvYufNkPkslYQD6p4A1OHMt5v9wZgP8BHjxkKRT76
RAqWjL3+lySxJGIiDXKtDh1Smst6uHkcEIYIS/B5roAerQcfzC3E5LDjvINqG6vccbOFdwETt48Y
CwYsmuRNfuhUOGl9lvQ60xjcgxU/zHf8tbabzmBAuSAvk92x2m43Zzn3k92khbRcFqoMhggYZKUr
EzXUedKZFg7OvRihnyRKt3wqt+Url11Vy5IO90dMVdTqzZ7T6TN4XIRMfzXSPXFhRVa8VjD+y8q1
3HyMIhnR3LPjuN5ujsGG0TnuWXWWhRttBlC6uQQay3gJW4rxcdzohtbOuJD4o2SiS+9dd1gNpetz
jQJWJBrU2V6NTR/92GKPFTHzOdyXdpDKAFh0wABfNj3acyOfymqzCc7C6MrYwtoIhrpHtVOVO2l0
gRAZYCQIFhIcETPeg/Vt0BEL/jCefnw6gCmQW7hiHgddj0BU0/j28JiQ1ib3DDPo1n0Sb0awwrHh
bKC61JtUx8/VBf28SYlhMqbqQuBS5pJyCxyOnVAxshzHw6fM+7F9PmCNE+eNvuDqiF580o+VbOR0
znw0UbI5BbpvBnsucbEdfXThFVijIOudkT8DadVSjek/qeJm/+EUOE7y+cK82axo587ISeBM3hZF
VQ/6GqSs8UshmXSn0HAqNv0Hj+ZFa/hbBMBVIJeUnNc8t89v7ZIeA0NouS8S/GkrYJN7cP39JcNa
kwh1ziy11iW6twJht/cPceZk0m4HdtcTK65hauAt8KXx5P1hOGFLc9gUbmvr8Gv0H5LaCfUt98tF
psPE+9laOiPZrNL1jjoC+qjt6e/j/ChVJfwiZ59DVJUv+1kV7HLtcKSJoyLR9AbKfbRXb18OySAg
ORizb++zKrk7frYwHzTPfuJEQQ1zlKsZ/yz3zA/MFtZ5pYzhrVK8ZarHrKPts3RFzVI78BKGd1x6
I1A2qSkqyq/0jpvNVYmm6w4jwV77X4eL6qVrh/FSyFmZzuMuWPuLnWQ3hMlXNqrl31rHK0pLcKuE
ILyIELRiiCxC9jEYQ6TZuN60QOrpsBkcz1kjratfUCGzgNGbcjlZCO9i7tRzkWOvu4VpKEwfyYxw
CcRwSFdIK30oQ37ESegXVwPJZInW4IcL57/sLvN5pYs+m6Zr1rjwa/ix+CUYEzHC4cF21A+bcn1m
v5clb/Fc+PvidKY3LTpDV+tP0qN5rXKItt3mVEfRqEOHN8dFtu/k/aJdW7ybi5RlAsKwHZ4o9l8S
GTijelW3CxRLd+/0fi+g/ZwQ5M97bg/MtZAHdO/AWv5kSkMaw2SH4xRmBA18KlV0ssTwuItEPYaE
RG4OOLW2pRzZgpi6M2ody+Ya+HqkuMN+e+b5yFGXfpslzhZWssr/y4MVRIuEpdD7Unah57iXTr9H
yNtjOdFG6tF3pZTokpIIkVoZ19m3GvOTDOV3CkHifxZJY63tZNfkKgzSTavgMpB6MXBTCVvxOhwT
8NIyPpzIJ+HfT1eYrC1SCI73FUiiE8qnApHGeQMDXlygRXgEDBKVEYzJq61FOSrLWgDyhTxJUme7
Z9oia4nufuQUaVghFqq45NqHS2tbrBp+BngkjmEimTUTt7jgtjzSaLIXR1a/NdHc4VdggyJVg1im
BsBV1K2phOKrCRNSMzWljEVbVkSxCJOFKHbJkD1YTJLNzOk9qyaiBWlssk8akWgm8TVKNmrqtg0j
XJdI28qfSdICC5mtPxI7OCPuLhMih00Xbb7kKLHIxVe1YSzjVp5QAuJkQVoccdjrIAUdjxZNhxjG
Fw6AmD74nMFZ/7b9gXVy2mV0esmS/HA9sknHqrgu16EkJgOp3KiOkpp0qDL1bIF5u12IMcbcjp92
EblP2pJsyqrIf8Pw7afF2zVLMuJa4gdT2lWqDItl/Ci1HKSF0Y3nQVSZU/e2dtZZ7dfIZDxdnQ3C
Nh8kDAtwDJQYqRTJP5fm2uYgqalCmzw+5rgkGEdvT/b7iAgtKxLpYLO4TClhviNJvF8gtl2aKqCt
JGxzxC3EFNKaPpKIFP3iFq1pRMdSQxaNyOvGq3Zn+uAfW4AARKkJwhKP2T0L1a/ZnpkNaXoZVj5i
4x1zCQbtumNCVD+/qtwazV4xaERie3GYMFWbIPE3ieK2q7iyon5+fpy2Oc0CX8xW4HyW/dxHkln9
l5y4aur0TazFpIATVL6Zm7OMKLMFYnAIti9oFBhYG0cQ3j01Bu1wNNyXP4qAG/+Qi9X652+vRGEA
UjoRgjvuNS9WjP0imAAfCk/CY1LnmBae0UefiP6b+3zFpWwlq5lom6Eg8Z2Ge6rSB2yxl4L9M+nN
6Y+g7w6JgUr+TEO4S6Ztf10EVcTnpT0s1Kzc4qWT9bTc5yDIAsJFatx+jbqe9CX1D2eO0X6qDlI/
p+hqwDBrP4gzU6TeOchn2kH2nid0ennjHZ70hOFPy1sIXpQ1h8LX2GxYyRA7A2KWrBAbBBesqtt3
ZqcQI3iNpqDNTrNlHPar59wgyDYWE8EhaWsQ26oZ466x2Qbqp1a7iJgUS4MEgQPeTeKhrOlqWr0p
UjTwZB6k26RtNBF4yWAktxglJydJO7aNRbX6ZuXV27+7unyFCVdjNooDOiiiIkvkoYeZuGqt/FsW
mV2msfCvHNdy9RdbS6cq08hPJ50qTB11e9avyvsYEv9DDBH/PMEXyIVb5n/2OEgpa4N5VsV7Jrtr
jCKaVW8GpnDZqQliJt86U9Pit82kiRqxJENbktm3oWIKN14ZsAVhg9/yUbXXsP14+P+9at/IqsSr
REkPARhLAOga2NBF1rj4Gx2euDfvUHAlOctnmbyBe7FXT8nYxGJTyDt2KqcRJ7xXYSEHo9DL67Yt
SSnW5VDcqN5oIiZygdVc0PVl9PY77Kx46lDqGcA6UhuXuPjZBcrpt5RV6TdxxNPT7IH7vx4bHQj2
+cjzh7TsW1FHJ9w6vQz97ADAv8zMZy33z5T6BbMh5VzL2GOwWgTQHiwp0u9DI5lZt8zUaJcMkBjJ
UGMCthuapHVbDULbBogvoeEXOfOcSJLFL4T9ik5ntbz+mDr0MktSNrWJfZD1DMvwszGkQHrizRZd
ddZtK4NNeTaJPhQHDD0mZA2835WJgka6clOQOANJ/1YTK2zfS/pUGAwnY+YaRzhUIXLQ/87FFDtM
106MtQgYGSqhMZ0iQugYCOuTvjqc5HjpLexIo9S7aQmZlmoiaRC02kJzsa+bm7VsfY0+3xLAfgI+
Mxcn0IhAoteJuqDlWSaVsUngPjLKr7Lo86VeVKaAt80fylD/y4nKz0GXnFaOrdHAxWQfcsu3lJhW
XQU8W3SYeEAunxoQJNp7Yrgg2SUzi4qLcKc+giWDgVbnj6Gr3UvjcN5ZzeP/8+w7E+qOWL4ifY7e
hJymG3cQ9pYGTDgdIq0Gz9ipDTuXZuebY6kWlU4xtjf0YSkpp+g3wHgYtDG8PuPiAQTGj57dtFFe
bcKcfTDMMkKhq1/xAlMg2vOb2h1SinhO4Zf/pnhBvKXNj4arAATvAtVMKlroguPyfOcjavUaLnNk
KhfxWKGHGDme6JR6smH82YT6y5PPwT5M2OakS8q/kPAUKdPfLbxGgtDTnrzhfWywXwV5J+UDnE1s
b/aA6ZVZtY3hJU7aqPO8YuixX1kXLYWiW0qVuNyUnaHi8CSEd7fmEIXBd14yMjwUrLpPcXUFVpek
iyjMTLO+7zXXAc30ITMgS2MB7bz/WxKZMrlNV1PddcexN/RQRuxmDKF54V0nazcv2ZNrxLvjbiNh
7vTD6LfvC0g8taC9aQmramyY8btoRGoITwVroTKsjLASwfyEhJeSEnehcEKqnmV3XI9yu5lLqyfV
pek7L/p7ZSnckn8snRk8NPFtx+cdACLFOF9REbS4J5H9wGFioYVikwtBBusKeoGIxhicgfkSqCNI
V7S75JgfEo34DiZt6PKbgsb52XziMJlsBFrcTpPhEEQlDS8fzx+qQrNgo1N8YOKRuzNKTodEGYF9
EibhmsfFVaYf5PRX1m/87u9gMFWcEKKvQUzDOP6Q+xplnteV5K0uENQ8NQ1sikDQIFdVtiRfcPhj
yOksz0c0VUxGgxZqmSO46wHFgta6U/bQUJpQiJ5yPN8w5byJtf+JAxyHi+F+UUPyjg5+rr9/6D2j
KrbH7FUXAs79l7xHbJP9GDaasHGRl1eAI0ilUTWJ397eza3zl3Y9rOmtmWZJpWsvt9U7tfpyMgFd
WeSeGhLZYJhcNx3K5LvaK6BCNQaTE/FxnR/NbJHqmPCxGAq0vjdebzjXwkBd5XY00l1UCxL+w0mF
VISGQfCWg8BP4eUQtdK11iIAhdxsOsZSrEaJS1P6kYK2rIYSykwR7bvdRH1N7qELauoKqNXDpiWE
cp1jyiviYAOS3Qo2eiglroTvVHe9jgUkv94KcNTB1ETfRD4q7N5WgU4m1diDm9Fs6EEDNi5Pb3fD
6kbpP/BKPJ6VFVmvc8pfRjPrwHOhbWH7mIgqQiJw5+/G1yHCcr2Y6MMjo3uFbzI43UFXrs29ABDJ
17mn0MypnKucmsBm2L+g7uq2pectKFSDJutF212ZJBQCRT6F3qC6YOPB06ta5o3NSBfrYZzBthlQ
ed02STPRnRD0gOKI0dWsXTt1uRRHTBak8OKXgbqoZEdz5yY6u7vtFH9/AkMp3oJoNTPjZ1sQ0R3W
KSdXx90RbejXv6QXenvcuSZrPcj7coWUgfK4V2oIHXJ9/Ky5dgFjsDWzgRLJAPtHYSZqlXzw3ap9
ltAXs7aTf1aZEYPGhcCiQECxqQ6m/vWC2QBvB9KH9bIYi4YLFvRDgrj7tevwJm0/GV0tUCB5Y3aZ
aCKKvx6AVa83rz+Dhj/1VrMHsICHZ4COLKymmaqxeBYRMWO7xszw92FSL5RA5NO009hbLSn7gmMe
oeQAfbuAso93thTh8oXN4f6PCdJV6wwtYIpiDM4b8QUj6E3UTH2u7xRTrjTtuVm0SiSz2l4DF1xi
Dd/p3WwXUbLQW6N1L39LGk2OoZsXnEf0g66sEatdiYgCIYldxjraw0LbJArLkLFufLy0UrH6QofZ
ntmtti7R6LHWzSxZ4ArjpCV854H2kl/djpg6XJJ3UO+D2IFyJFJfeLF9gxaHMGqiGm9rwfuysD5G
AUNwL+bOI+CCMCN2FK3bVTQmKg2+S+2pRWCNClwGmn9rTdPuXO/1swv6LcczQEHrYqR5EvRR4U85
qu69mZKcO71/LRAFmM/yZnh84FyDSfOJhnpCHqvTYg5neWGEJVGR/F8EKOQwQ70/QtQ2W0kOzk1B
AhIr2/2EIcRzj6DL5a162CpEvWJzz2WlpySQvpJ0fQCJ6S3WMEbeESFu4CoLAB3fW8L9HHhBjkAg
Q7HhZwsnApXgS+SIVDLLKIC8U3StdSQq0uSAJiSmakiHCObnXm7K5nv3C4M4WpDBK8lD2r9on9il
saYHheVon7m0YUqTpbc9yBg6TnhS+IRT9cL/2ShVbtwXWLeKes/f5KJPg2cMucY8pBGjNwOsyeWn
DC+snildTo2McDLo1XyGYEDdOPVvPDj1a4hX9Jnu78ocKSoJA5jFqNpZaujdKcgYQOHsPa6KpuZP
F2wHbCXpBAJjXH3kLFmt8ehCodqzYefXwB9siJC2ULNmJZ+uy7OU5zkScupeFsR6NmoFNlEWwsGH
WqnTUWKcMDY3L2KSJvjFuF0GylR4nrmBWELJnkOM0iF+uFXAv+lOoGyWrO21twbf51aI95P3si3g
BWhSJaKaSxEPKWw8UgLDeuop+CSKgCVViMa7sIh+jRcoCnTUhW+K80X0hVsYNh3G4HlwHz6yp65P
wAfu33HwX731YPMhBEwul+E+ARyuOYtrAMkymF2zHAfXv32acSUVh+cEE0L661LVzUPVRkqoebXg
3Q/rdedhQdhHm5JWNl7k3ShxeqokloXG8rKy15CQbmfouhydhHSeBHj2vu98+lNDmSZHUxThXsg+
kb2VvC8+QHpuRhw8Na2g20FSF2wGzb6l2mqa1HV7asyy21wrvPV8+ZPqHeNk315Lq7w1xOASacrg
WIKooXIbtwe4Pb4lEFoQIiO2nq0ulbFK0Zj/u48ftoUS7AaIQ7LX8SPRSH52Qkio3qntfR6+cIz1
+7LAldTxrJexepzTsmsL393XwHLc6tpH65I8hD1OkhKejiNtG18VqQ0yGF3Rt9vFwzJp1UuVCfUx
00IQXFx6h+D7IMPfJIxb20K/ljdi0wmTcI/Q22bK+4PZpyxJCtJDPIAFG/9ZlbQ+UDy8wxiJIBZ0
NwPGeFVWEAaO+6yjsOHyuhiFYlLGvwnMA0ueMFQ4r6tnNQLR38ozBp0FJ/Qa42HQKBv2qpEg5kRd
Ku608JfY+eqJTcTV6B1I7nMUbWj32APTlxvLLL8MgE7JiKt3e+yXpQu+4gr8KUHoUww3IYAX7Gdh
5/gciSw6AVmLta1lZ5ltbCWoYsijk3RzKjKdbBFpmYRRBEEMkaLHsmfuF9xHn0kSzkQ8eLPwJA3s
XSxG8ozrJ+jequ4eRZ5CzgAWpO4vsB9e+CzUvVQAAVBnBnkHmefQzPZ3ySAKbG39jldlKkZHLGrk
7KBvY2V+oAjOcjyvh35ecAKkJSgI5eo+WEFb1PpYSL0YbzK8KmIQAMe4RHtKzSD+/BxFJzZ7q1X4
EWLZ+kz8ivfUdIWDhuha5PZoV6IElr5OZ5laLREw9nYKhWRI5/qrQf/H3qwO/N6T3QFWbmvCmHol
OYJm/KdtOioOSqkza+5GVxK6mD16itjXoXkdXh6Oe9rdlwj2Gr5e8BwVFRooMXaxNPG6YWLXBO91
8rrlzr1J5qkWO15QGDONxMCrw4M6VBufT8NMJf+JiiarAyQODKbVF4Q6795a/yHCi9tXCDR+8VQz
lF9fqpruoeypmITU1Eh6m1CJ/y7ekqRd0cK7k4H9iDvadTZzdM7FMMA7GTe9ca8FZm9CNm/Nm9+S
sNRcoDxHu/4UdPpDvigzso6whbVskn0jIOQvsCkWKQ9EgxedeLff/+QVmh+uwj7LpvOZY9z46gbv
X+pZe+JmGWvq+u1yKhC1misjNn7mr25pnGElNlO4wawMa3el6sAaDlYXKFVaBLEuPRMyfCcjvfNF
fYlnlweoeUqRpVL+rwlFW7dXgnIL842fX2UENQboVhl4Zhge/L7O4jmHrIvYCihPuz4x60A3tSYa
Sy7qhjkfGPeSn9bLRujchI3irrzNh/GRDEgfjTGYy9ZqCc+SBFv11WC/PYu1SZJTV9atiVf0N6sj
VUDYhSgEQ9QqnO6aadCFG0rTOkOR9yJfLeJeIqDMWwURW2sYJE6oFwsJB8GuOhmUoafuLBGWLe9v
OK1ltb3GC+zL5kZOXRprDs/BNiEeSa+NCflKMCXGmfrx9g+nDSkP2kEntWMpkPM670uFBsA5W7V6
2NIPmFfc1T3PqR4J4uyJ7zqXxp2GHvj7WvQJc5yTBVHFGUkI+9/RqLQT/4z01rgDgDshnO9dVQx7
LBhG6ACJljuq6H0q0phUEqxr4+4oo7CyOk6KV+3TjllGdF6urGBTQ94MwHfeIf3xhZrTBvMPVF14
bjHZwRqYZpWEozCzQvRP6UDChOlWO79y1PEfiui+JaLbee0NgA3XmE0yDXBIwn6QrTxCTMMmikla
Ice1LyX6imSyfhzMC/Yu4yDQdskMghU8IAqzNsQFtNNghfgFu1KCyuRGiqUXaeOSTrXlPwvXzBaQ
0B4flmZlQiRP7ho2npf9Z9OhpZwP9Y6wCu3R9iop7iZSZjvoWGpC9G6sPNUZuDdw91ujhB07kqG2
7juk8Lj0hIclwdNly58Dhy9EUkcg8Ul6K+Q4Be5fz/G8l8diP8IPZ1qMaoZ8fTHfbvBM678iW/pm
ndf121a66cOYR4pc8Gf8n/zbFpEueVqcmmLT4K04/jOe6d9Ef+0nua20eJRSsxbdYzYoBiKGBbQr
c8WxZdFubRGjJqK5yR4puzEiix7nb62ynW+svgnCaa6BeODlL3J2qqEzJcJyXlqV3fQ8md22mJmX
59h/xHeKEhtUVms6U+RvQhx1pxqHQVIaItrDQiKmXzEBiCeD8vGjIWH9wbpj0DKRACLf40NDRLqo
lcdV1DnAuHd0KkawqWixF8dw0ugNTzhTKGJhKnoVMMIBmCZdD0Iz9ovHRaOFzbpl5f+jbRP2bjyf
ba3LJGG9N13AL8Ln5A4vEdsbqtaI8uVZ7NQn5CRIUXYst2e66J1Z4fkTLi/bZobsQGvXRYm02t2V
lZD+74zUGOiQ8GF+TKaieLuNQVaYNyrPPZL+3RwhqztPkMrT6E2ByXYVerpmgb9YG3UaoTi2HXey
T/T0x52nbvWgCwEsn/YRGBNXllCTMqPjoguSAcivpW1rAbnRe+b/Tt0j/AeYtHIgJxlxMgWxTt+r
NaJ/EHsfVmOfi+V1ecZuHNd7CDGdJ9rMdhTmRAWm8hMMAvQL3bvk7Utn/jZRHOBksvW7vIofv6+b
7FpLqiy86lqkjWlR7pjclK6+XUzA1CqJR2z2g+s2fDcXv3T9U8RzeOngijdlHknrSP8dRIEkesY6
tJbDncjta+0/zkyTYG3Kwqh7aqOqYqaCo3AT8+AKXPCgf+uc+ozh3/Xjn5YsgqWDIcSP2WyJ0L+h
7gsxduDRwz58EgkOmjMZth7KH6LMsDuiJZwOvyzxvhpUZa3gTamZ/mCo9zsOGkX2iFTB3lHcXIRf
Nql6EDrUjClUxoYXZuKhmwMD5zC5d7dl4Oc1MUvLZZ0NXasBbyRIBLjBr6Y1IzBTVpufTszOjHOw
m5r5LiXGEJ2CY18YCjNXgMfhZLsoHPH34XkSC7DYQirKrqS0/MZy/CVQ8LiSBqqd0e/xtDaM9hBS
fQLR9cqlyEyqrxp60cycNxfjfJ+GstGr0NKGE2xcc8e+jed1Hh7f41wgMlomHw1jAJMqeSYg1vL5
U22MTyW4YZ4lBmsmkmYA/GOBbgmJ3j5q1VkhwL5q+SSA1+/xNFjCxjECvn7xt6WP9qmsu/mvUCU8
7enz9W73sOmf2OpEvyo6QrbPiRES9XwAFlvVXxGczo2dXjzwCi0BVCe/E+18/GGMc8QokmjTDeIi
eu9EYGt2i+qumKhwPaxVtQNbH05vBOrBmTX5dJ4pwBHg5UMAlczAEOlWbK+IAH1xjvKE+EW8p5Hr
9aFKUYE1jMtXgJYXTjKonSKBn+6pcK3wWoffD4iDN9QPjd3SfCArRgt/FxqIqmbv62oH+8hELK9c
q+4ZpLxg27M9OqkR3DNsnXtHZMiU6PJWOed0lZW9BXk8W093LLwevzLRKZGuzSe175Ugg9ECM8qy
f6QIyMsPl1wfspXk+EMVix0L8/8vonggjvUtapiDrJTqWE9nLxC8jpEVSGRURWQ/PEqbohhC4guz
rq7m6MrQFDBgLPx7uR00tFH+at2Owe2xBIFD1NC9tDdcr9L5lk+zlUUnl8n0M8aEz1jFHD+/12lz
rnhE6yS28mR+f99F6pGjcVejDiW/nQNVnKQ0F7o05s5HVZPcYz4z+GuLxhsKBkXNSQLf2eUSDMDn
+0j5HbtbZKl7sSs0BoSbD1D7aP6NuBjFcIf+84yKALqVXvyXXiHlYoaB7YtIIir69NaYsH6pW76Z
j3CPkMqYsL4+xoDe1RYOv8oPPFFrGgwoqCEtwnUkIAlmLTjXIJCaK757p3GL/B/IFhRKbG1PXStj
L0UGSCwTE3M65u+LBozwkghY2xbFoxiClfAey0TtELQ4FfJc+Pt1xiDozlgFkdqEy+aaY/V9hJFr
0R8ZptowSPrxzkm9I+ydcBhQuPzFi4k7lmqIX+LLOEqAUWW6T73NGA2Orf+EjbZklXaAcOfPF2te
zqLajZilHfbn02YQJ66e9Yq770fdjdqXhowqV5GJKkh/TorT4NmuIPhPRvnm66GS56cDp7UI1upS
xtYOsQEik2xPTttGzBT6BPKA0wjQ5TbNt4ORu0H5nwmt/mjS+juYsDXKhQys0QadMhE4yJ/nUw11
vQGFLFVOPCMrYV5Q6ONoy/8qJPzWY21ySoSI9jqeqfpAVFjUeE9AU99QgsS7KUJ4KV7d1K1j3X5Z
Im68EqFke2piT5wnsuM97ZTnaMVH/3hp8xWMYRl/LHbEN9+m5mEWUTSZt8c+knGQ67xxGkl9BINY
lOH6hJ0DwYWCuHsigsCjGHsRUzt5SdyCe6EYlWmpituOqywdzRP62eHQ26ih1GbTfYpgHTAImO2n
tR1uel8Wl4ltkjoJBYnEcMTxVUb/UKODmOF3U1NOxbYUBXKlvpkgJyYyAx/iDp4ByQueVkE7ZsWq
SUVhLw/ZxmTn1FrJ3VXLgjhFNkVjlmO3wQdTtsImdQPu8PGj9ahzcIf0JG08XHjOB4kLUhZlRpRd
iS410dzz+7I6JIdLpKv5sOBCmlC/k440YBA9/X3ub0ZZux6VRcY9ZRsLAWQScavNn7WGtHUWInbC
XtUHJ4dzLfuZkXUP863dZeC932YPoJhyL/yvmKNMVDene5Wd4gUaerK0FHAgBmGaN3XqaXpou3ql
nZJb0E0BrcDpLEmCXbKif1mDFyI4nmgQ+GVdrEbNL/x8btxaEtsHtg4ofwqAKng0wV/79QdfhJya
wFzcNOtnYHKYyi5QDi420aW2DRUtc1Id6CZBM/DfMuXLgLNQFH8L5OOv+6tRzoQRvBJl9/po2ncZ
rpSHo/hPiWr7wUBc7Eybq3EsOWhOdjo3oioSR8qxSdjAV8nihYJRWADy6D+hTPtEV4XaFA8yKY39
6KpYv6Ix5RJzYGtCIhFM8hwHqTbbdmBZPP3PUrxsY/WNeaFUXBaWS+/RWiSmF5qquM+WqesaA5jd
d1erMTEm8ntkLtcC2MwRtZp822iNMOq8w+65K7ZfE2PZwmCRCFjgjk6Op1Y9HNSGQSs4lfAvTNOR
DfMbA7LxRHwXPWc+Ba8wqCMaYZhLLThUSPpXTaA2dYEnOd896Md79KUXkc03U3LVsB3vqIOuvt2N
swVtTyLpUfQvc7ljY5E6HC3AdtiOSKnvX27rEOHUz2hgxdYk6t/i0XyxkbQ1H/f538iq66hFEGus
6fxhD/vUW8H4lXnSIaT5HaUhii+RhQrhC3u0567YapyhobSjXjsUWTN9Lt14NYf1Ygex7IHcAF/c
UxZy8UQKHu21T9jgqHfbfx6P37TA077O09tvUK02Ika9EMPO7qNb/KwiGTeZgXGC24I9j/DOF8dW
OSjGUB4sYbMhimD08WQZR1NxKt7GHhiDKqo3KoU50A8yBOLLDiVcii+kvuoI72QahcpA+ptKpemN
WKjJ6yYQimtfzvXPPNQ/v7IwiJ6jx0fKRIhcSXRhlABtuK7oHkWF9HVVnKPBCHQohOl1nHQEdxhf
x3ugNK6KQbMAFThxX9EAydoxFO3wpxHfrLcMAC3b0VaLanTeBvdOZSq29FHtXyDxzEuHq6CcnWFL
d4rdFY7aTLpSMXvgidWOEjtoIgpqzonS1PwM49taCqD0suswYvnLU6jubHpwszSlVX9A6onjPJeh
Ws3IqurqK+DExVnz+kT4ReMR5gDo4MmkabJzpR6821HiWJO0xqsi6EaMivXIAJ+qh07Zz3kBrmtz
MK3qXaDsxaGeFsvKgIxF0If8Nk6mi2SlRp2q/pwLf0UH0TA6qbpBbjF/dpZwUZlZeKPGrpjxLQey
I4j9/UcSM8TLkMgi8w/vt0hOm2+O2bSxnJF8jyCJfEPaayKptBbavfzZvNlO4o25OQLx/t/wMT/R
HyGXnJNHdH6cPDRfXBJpBlZ8/2dyPnaZ0IqML+RCbYw5gMWY7RqmggWX4hDYTnxJDkKiloybIUMK
By7foQEa+EfCy1gsK5PI9RvYa96IcKmlMTcCkwWiQcNp06drC/J32JvbJmPAY+uBFwOLCDjSCOsu
LXzOkJiOQFFOH6buSU+Ki1m6YLMPs8akZFz2rHEfO1qVQfC3nitC88oNcfzjWeGElIELEM3o6Ntc
PfTJ8hfCn7nu8LeZm6116QgGakoS8qDieL7lvkRNupy5/3zxLb0gzjHC8UXecEvtkcAYt1gnzBjH
GWWtpEAtKTcBjcJjlOxMJtR5JYEEn0aHOJN5w3g8vNoHN8RFVeqwjzA/N8Pklu5fGB9HBMp3/PmQ
kIdkPrODQEeyT8IsfQnY9dJ1QQMRIccel5351jl4L4kp8J6U+GZtIK2SfqnHJKQrsyVbTvRPvx7d
jPdklbcZQrrlZjbNdB+doqFeqNdQxkWkvrXP3ekDcPgthljQcWIG7xMl8EsDf6zkXIzfjVbigY7y
/FCOtHXL7otDtVUP5htQAYOJcJuMkiB/pdDiivXHxNLYIxEcXUkp1bSiQW9Jn0rSqx4In66seU4/
7XNxCru3pm0dMCrd4inhc0RM2h5ovTOx/W1gqtwwOmbAYzLn5CdP5Zc0BT9Hk9IP/+XOsvPnKK9a
Rlpst6CpM64dzapzNZhKATZz+NVDQf1dOHmGE8KCDeN1BvJtul9W4qhfhABbnptEk7PTq1QJZj0V
SisLp9WI6j0nlMw7dyetudHavuIRQ6T8IX4VEWdUNL5JX7Z4Nuzo//pQRWznUs5//6K/cCw+b+/7
LEQERAx/fvoB38DQcuf9Ix+5dxy2jduwbcN35eJp67RjvN5KwxjNiIRICjfWEarND1jCDaZoASDT
RyRb0wxyA7g/g+MgyZBoEY8yvTpH6J3mSME6rV7A7b3yNOCPXJWNDFIOfm+dU8K4Py4Eu8rQWohI
LapxaonZtERt2QDEg0Rrm5bYfvDon56T1PKvGy3x2m4uR7YdtXGE95a8nPDEgVibd5RpU/I0lwWZ
HufVClXLGVESjrspkGuYpP0SGMCkjfZNRZNIx+Qr+8KJFDHnkeNVDr45OBPqcBA8MMzBDHVomc43
dlYOofFUVvWfbkJqMKGugEW1hf22ANfeNQwCo9xl4Ksxgu295qWhzsBZMDLrIbIzBEhP7RzRbPhM
ZXMo2q4Yol+q0L4MT9eF3jo1f22c3XYSU/modeBtIoYupGKnv4JgDiSgzgXrLV8Z0DnrbpYZGq3m
pNA+RE8lMgLJJ+1cZvMwaY1aK8H6JN2wJfArlbbbEubKKp9JVaLsnf4n2XzPnxqdoBMDtU9dJ0wn
jm0jCQDj+H8APZGprJ3Sl2ZFW4g5nhkJupQtBHOtclU/F3t4eKmkBjdEki821C4oczfQ4TJsKJpL
g8XNiGikdRKsygFmKhpBKux2xmeFbTMtJJtXX008m9adiR65RLsP0s10b9Dh3PM6pa9pVxaBnWfT
JLU8++wkGkNtn9PxghCK0VGAotys5pXrNoP0an2vklJA609O3ikFtk8aPEYBJfHcNeLqW/M5aEYO
+5oMR5kJ2JRiLCfhpqCRzESupCm1gyjpjDNe3++iI/J4C7R+asEoekx1m8//dq1ODcUMzjW+UPPt
/U5kvFKE4/7hNWOyRebURV9lCJEIG7H14K+5SOeKziBfcvmhEi5svyvEB6z1odl0KwAC1+odalmy
ItI3wcNRCRqZzNKDmh8CDuAKHFKJ/ZIoZLNnlNev+v3oNKaAyLY1U+hIMoGol3MtfdWb9vkb8cqP
CSh7AlXm61IxR89MxoqktUBkBUwO/v4xlJiO3qgMLyGQf14sFXH6VWOKTpX8c1h0v+DuW8YXyibU
pJO9MCu23QX+VEAwYV8Ls8SnmTsjMFPnLb4RJ9VhXJggLTJn1rr8ZD8pAl1iH+5NyA+3z0sLvIG9
ZGxRb4c3eSwYFm/Q9KiutYPlfew24cCzP21X6DGsZDKKAca07N7/4ADrkVC9zyIMwbjJhuLQ7OPD
Mc6Z13CNTXzF/myE72hQuAo6ireZmukFSc3eVDX6RCdn3UtSWXcWU+9Jzfcf/zXiVW0E/HfIHH7H
fMLj48DCe20vUOUSezHGmYKCe1zwWWHkCQ3efk7FLeYluM5+c/qdwLY5JOMtnivYO8GwO7CWA9zL
e+1MhPEhNMyg1HuNq8kJ8v5f028Pz8TaI5aIvQEa3qdB+3tDnezbzPcQvYR8cSu3203/wjrAD4H9
0bYxctyz1hxnm1YcUSmodXhzHM0ge1cbR/LvKIqVMJlzG8DnW/ZKKdDetfHPJ+T2JzV0gbfDN4mZ
Kxtpu6fQ7D0PN47RMWs4Reb507Y5gwQeFPCIyNujdDUuxCnZW5O6Czojozt21mVmVRRdGIpIQOLO
OneKK+gEZKu/xkSMFHQjRRy4kO02zPT14WFDTJ2LfyZjGraspm+rFpczCuGlBELjkLUmnKqfUeKS
BMPhp81bIPbJeNlnrbWWrh8ILAwC2ZAvnfQc+ZWEyRtX1kVGljYPVbrrDiMBA9p0madkH56+XfT3
DQ21NkyXGskexrlRE8jWLZFZgFh+n/iRKlmGtkNGJij3k8wlPcwZ4alNYovnoYUuLFDLifBK9wq6
QSUEGP2RkcPMzfjLw7nSZ8dM0qohzeZcaww/GKAxAvVaq85evlGtcP5/N8JmnBavaL92nzisSxkW
5WSPs/cXcOXE+4Hf8E7BPZtemGCLLBUBUAudGG5DyRqKwT2cIpg05lqbnhq4T4yFiQoPCLdZ1vMI
zENFsxp8vQanDjpO8caQLE0HJl1KBlN8MNomvoDysmbNmg1Nrsoxb3uqmnRGPw0Tg686TM1548WH
Ua/izBKAlLE3Up70zZuRb7NcCwup01QLFb1SBrrLahhW/OJ70EVGysi3RzYKF1lRxKNAPv7Y3yUC
v5qnzRcoFAQmrTQkr34s3GydgT+nMicjKouHMUbiFNEtgP0iRDLEJ5dwZVnzgMY2pziSBql4T+b9
RhJz9O+SKXeVEvIJIIHvr1ejlVRs6JJ3wG/KkdYG5NbvPIsv4Q7HDEzrw9wu87GndrPGl32DhejT
BeF+xi/I4OkUVihEJ0EM4JzUqTKifIZvzwVFXIZbOmIRwVFWspfeGV+JjV6LIyFNAQgHHB65Eif8
QNbVIuagpCXXOyehpd9fbIRs0/NWvjMkmp6OecRl2VQb/aKz6nv9mO4JZUE0rnYR7VUmlz6EJEU7
T50huxeYsBpYRVEs8zpzCzA9276K2IobPcJtWFLSD3RxXu3dvVk32pPqPBPSb+FGn4l7Ep2O4Y81
722dktaJexbl1uNAgeFsmDcjM8DhKpmpifDXGK1wnOD6tFaC4mfFpv6YT3EDNFNJh+TCPfQ0q+vX
CcABCgRKMRX3tiW8u3TsPYippDxJ45MfumSd/lj2mcPtyDbY1ztfFgkFh05+/dYaTHIWgcMpuIgr
8v9726LLdTspYWUDOSaCF5VF7chSYpeadla3mxD+crVIBw9Ot60ap3/ket8br9lHtMAPACp4cQIv
7YGVEXniZkCDvDABnIlOVKrPSMuplwhElmRmHC9Xl+8PBXya1eCXxORMg8zjmlYbKSV6NMkpW6dd
ReeUJADQX+guiw3HTKIQmqNp+J1g9QZsvBIXq245dlq8zwYXZtyNadr1dm4oo/tBGYaVNnZBT7Te
ZZt0Fa1HGQ6JxdW5EHxvN0Yx3cX6QRaZqEgYMCpwGiDeox6lNgHlVlXmRMpN0FdSpwN8sCDNjwb7
Pjl6HPZFynAz/X/U0zxdc2o1q4EX5px1wOmpJBYArMbH1Cj5VKbaQcVNg6gvTz/l/PWtFfmhB7fV
VIPTrifyIykjhFE4rsIf/TXWKcMcPiINdXfioJwzpU4LvKDZztuEbnDJSRWsJAfFC65zc03rwdC7
RZNy5zLnykpZKT2rRazA9a26N9yUnTwEh4AMV4xZfff7E33K6FMVwCJrsmaqmd8nPjrNvSC6gKg0
QHysRvHN2iiNYfiV6+rhXbHesxjwQjEU8e6HR1Sc0u/30R0kIl8fqblK53uXGMvsPABwpMoxQliT
7rnJabv3r8gXDUOPEr4mChMAeF99dNKYPM8IXTmMLEXgDOX4wr4CcueJaxI9u+Nq0+XgZXFTuH2G
VzwRKoCJRRDSUN1eZDMuNdVyN5dUg1b/zRhJbSIU4R7cXxSzctNlLGr2/tF0mvUgrkVRvNR6GOSv
dnztIOadYXBlioTECdT/UY3Ifdfqq3k3veBaOuCYKaJj9FqFWDE2nAjxILMpeu/g1bVRcn4rAvLC
avD10f0PiSpHIRoaZkD1QW2LWSnVpTWRd4XMQGp2f0yitH9OPh7f2d3qyFTAkRN01XsETzsMn+LG
JzIyKlWDcJWWBqPhxY5iE+y5MY8WeiGqzoJnaqJgBTzdH71ST0feLA2i4h4Odn5MxqUscZ15MOBE
39jI6TlglFVQFX+sNoA5uRXy94mp/k2qW9lA+rl7aHi/Y4vXW0uLRq5iX1j9+JIsrenHVx0+nL4h
Fh+TKVk7dMq6AhAU64aNt0pJ5fEV4W2g0WkmHiPBriQGCLmVPPJFwR5n+O8VFp3trTDgy+wntWo2
OKOXvrV2QDVot+A1HP3R9lMIxPd7DjXZLqDZqIyDm4968JuTHeoh4uClHCtHW24X3+FREQooA5GM
faS3fkEH7jWQOuMcsQaHogcFtcr/+FaZKEz9HdjCE0+mFSlzDZqthnE2sCCbKJYOgRLMSVbtEIGI
vjSw4YFtUfIRqFVA7eOQrGB36FaCoEOu2xcCOsBe1/Sm+gcKeK6S4d1WGszxotXkESWM6HtCzdSD
TZBkb8Zjn8K6j5h25+GZhlWFJ7Z/LRucJlIKOcMjPb9EQFbjmikpQtNjxzP9aW405UW+TnrEuKML
KKxb1Tl4TfHE8qiVC2Nt/+MtWFM5Wbbb4NvTEVoQU5qH7ek5vwRBHFy0SIohB6NDC6pATa4K0TwK
GRfu8iPQmWIVh4BlTsMNm28I9XPwdz+pxJVXWGyvhQ6bQtR3yHU0zdDuSQNPsPJod34xlgjS254H
d7Z2tFAn/s6PQmrw/vPoRVGWKL67Nq6AM89EbZ1w+gUuwGnHxZx3oM+eByDu0gkWC2Kl35bHEoQa
c0POR18+z+kE8+nxMTbqwqKjI2MET8AF0kiMl3sm37vQnZS40uYWkoUW+jr21t2AkRKuAkwAO4BP
W2NYItG/30ZT0DEgBdNMq3GgnISIrUaoE7H14o+93MtVCsrhDB9KTX/gT+VbndKu5HUufDR5kYcL
Fq52ALcHlIQy8MF51PC0D9zV+vAcQI2DGklMnQ1sJmeUkSeK53mGVJvKlv0TzFoVqE5up7P42xj8
pDXiSqKMX0dS7e9ctwj697EgWLluHcagrzoulJZhx2jCZ2hUkbg3n+wq5bEjwrdST4Zi8FZbqjvs
cRFoFbElDu8hbCoBLhPrCQ2bXmzeftfGeL3yC8At0LzHfLkGlqRVbGpyb+CY3+7Uk0674MCujdfR
rAuXAnvPLvogtPSKrYLHMprgk3IsjnFFQJHhwyWlQ0qcaimqp5j9fcY8VsHavXmYGDIixTYCjnKz
u7/4Uh9L6kZV+XxGuZUcrpmZHLAxoDZl20UIgj6a8UZKHrpspiInQwyeWvGmldwkQ4ukd8LCkPIA
mVPQrQTIa1pfYWQaWuxkC+K0x6+pdh7fjVZP4acnyOie1RvWylOIHOheRgtMvrvqQgdKBewM48ZP
D1XU6lgj2eI03fNL4BfqMb6fIzrNcyGvx1MM0LHVZxnZu5JDh6emz+b6zBXa2y03fJwvo26vWNEC
jl33xpl4ddoGQu+L7aGS4Lq0imQkpbsNIRRpAK0dYnj/uUa6rnbOxKslV0fem0vCErtMmmlvoQsr
IA/Jj2M/Mcewm22b1XBiVwRCfFn0i/0tb/s5EnmZhShv8PyplrrhF8URc5WNPDofnXu8e8BmMvdl
sW8/Rrlc7aYhvwYw0uNrCDEIx3hcSLe4DphlXs/amWC6l8m56sxF8/9GKBQyZwqrqRpbw8vVikvR
TV4uR9kZ11aW4eJFWOhepnlAG+bCm2ccl1R5gWmDX0R34iLLmt/mLjSkCkIjBuB1HXuTca3F0XPo
YwI08dET9Bd0JGq8Wb7Fwez/PcEni/L86bYq1Tx9eyGAkpu7oSuthY4R3bXvlNmKBBkFHV0OeYVd
DBcdH1BGAKWdTF5DUJHgBmZUqy6BR0MbzhhyReVUPqNTvT+5uDvGNNNqbY98lQIxWvNTkiOS+4aS
rHdLDnrkTUK4ZeNrItu7QCPFIXsoC8KztR0VE/WR5zxCwCLONIefDdqipxvlDqQMmhjISSo3X7yw
9nHv0r7X1R+2rG9HOw24vd9QwpjkhQWbBQkMYs0eDn+7QNH1v3SjzRSOWnu6DJOOg/iVRHuJkZ5N
C8czchsYPFvD9YpUfFn+9bBMvZNwjVaxHdY+emh0dynLUqMqDcnoNv6BoRvnqo6XD4Yr66H/b+0g
F9eV1jAwhXrMsrZe2UJK4e6Jn3nWSDf88V5vZdZQr9wr+KhYy/zLrqS6Jc1sS6cKxBy6abYrZYiu
pNoWUxVW2tT7zyq7Nehjd2d5uTekLvgrFIfm5VZMbwuYvYbj39wJ0y8lKjO6ykFE+5bt1TuV+3kR
0EDF2ocvbX6fwX8bMbllP4MmmQLLRp/LrpxCYkdkHqyKflV1AkU1XXrDKmyTJBsVYYyJ/W7PkTiQ
LJGcXq9EFrlsYXgSxtNxC8fK+bc3kCYkUj84Sd59D7tly0iWRbXs0l4RQPhgX5uNLGDUBQ75hHN8
Z7NdWX1r8w43SdFNajmSCFAebZpR9N7L/bXiO1s9N8KKviJ3Rwe6ovGZxJvtIT3qePNj9ysHJFCF
XSEFhZLgKTCg/9dJKWJocQs5DpNWElJbMpJzCNQnTNA/bTnXKELkjv3SCZEWxLFSwE9UXf6p6ZkB
HjV6gNRlal+SgBz+MJIt7wP7xGviE8QNK8QVCGPqVn3GT+ylezpzgm3NtRGPC4r6inxTFhk94aUL
XFHPZ5kMkcUlqqfc5uQa9RbN3XoG/VPQjtU+hH+l/JB7sVvvcbdiNHTEceT0u8VMN4zu40wsMm9V
fB732pWNeJNLLeAPly1F8IczBQpZDarP0lk37Hsm+C9DHqYw2AvAybezsQDHu3zIo5Ayy5t2oEFm
j2TWVDDNt1Gn2tFK/T+qdh8OBIqxlR4m+pgy8Zc82M1uiPTKImAcvzOJaDnpx/SuzFP5HthsArs5
EATFXl5ZU6khMRAzWtmaNATkLd9MuwTB2St67gREU7uiI1fThkFyBLq1surYG0tI6UorEsRjB7jI
pTWlXnaoaXaJm5pHtWFNXio9gGBSCDroPz0MimxyDhI8YS2b4XmW8CIRiCXC1ipSeGMBJL8jmDET
fLJnHmGa8tREa/IrK7gK2TUaCOLtCA2G0Idy+U7iRKrpiIpiQmdqud4QClfMeTzMSDMDdRwAZcrV
xbHmnCwU8pgJD50EauSl7LvyBiinBlAjDPfNtzW50X/K64K4xTE3wPG+TjUPJbfcWZ13cVbcOU4+
jjDdzk4HyA54XqeLA8ij0xK72ymZOaSs/oN60KVfvHhxytWmCMvV0VNk3kwvhoB8YNuBQqaYFr+y
LT3T9RNGPdD5caGKLhIWsOUDspbtZD234VxWCCl1+9k/XhH9pcCC/sBxdoYZyTdJAHpNxiT9Ok7k
vMVNXvqCicpGr4Dpzx2Tbww/AtzXCxNHYnaQYakcqtXfqWRle4A8D8n/xNDQumiWL4YzT9w+0Bhb
4DC5ZrtXyt+bpvtMdo6cxXxo55VxvxCg8cIeLtpwdpLn5ZdHn6VQbeXaf4uEqasDg/u9oLLrSxN8
1CQiG9v7cGOMfJB2o5lWA4GHK6bWM/wHSp6DhSk+EuR45OawZxDEsQmqbAoga9yhLMm/BJrIr80y
WLW90obS2ZFZ4cKE4EQoMl334XtelcgH3JeJ73/Wjvo54DISFjkyToPkoODEbg1ZDmuUfRSXBwy2
SK5FO7vfh9Zc+YTCx7zBDfA5PPXf2p5jZcUy8Vl13QV3elBw+dtq56+eXeUi+NqOt16UFiRDo1bo
0EI7HZ7jiIFOgxA9UrDRNkNurZZp4DGyFZq2u0ChJX1hDO+1AoNTYP2DsJ428nuQYWuRoKDjy7Ho
Zf1s3XGy5bJEptJ/3xPild1Z9NDiJAUMEeIxuWPr1Ina7WmIKp5N7pZl70INnnR0USypD8F5rVUx
MmfL8h5AaGCSge2YRFSEKbjJXwECrO1bWKiaxj+oZBGYw356UwXfBny3GyKu2dgJRkfJDhQvtaXl
D7gMpIa8GURu75yPU6twtqIDwS4CCZLVOpLRLlWHzRsBbepsB7tuNhovRVzinb5s2QkfjUn8vMJM
P9A9NfP+yfxgk5QUuTHTFiPLA0yc38PzWoGpEJranlpZgDua4bs0AFI0PGuS1xP6e/ThhC92I++o
SiiLDmGAowV4iV8DYvGdWrftzlSWr4rPDy2DmTJZULqbRrB0iSfojeOmlwknVjsNh5TRK/v17mOS
Wc+NgY5G4FZ6quU7c1VAPsc0Yq17WYf3+ned9PUFU2ss6nxgkMfBYp46YRh1zxiEeNf36sZ0onGx
i0Y4K12c5/7NsMGyeT1KVOEF7/vCYw/t8Kw19hbioEHVGKHZttO08KHph9sox4773pnY3W6Su+DC
ALYEPyMMYeXgjxTkww8+UqYG7j0TpH+lMmjICWI7RKZ76p0TRiD+PprG8ET5ppIlMeqWSIHEWhBK
dE5csxhc7cKxwm8XHml17A/d3NMZ5kaUWLDvhZ9rzQrdi1CtQM297jX9aENwdUsDQh9KleE8TYLd
tMMtDpGMRVL88hytuKWybcxjm1V6lmRG3K4DMHB2upC76EuZRMaSBQVSEKF4+jqNaNrtXmEBKkhb
Gl4BNaqOjcRF/qI0/xBd6z1FtJyElysS7wkFizlxzs6YYDPtZhcaECP3wkuwxdaCu3vD8yR9Vf1q
kwLCWHIORCufvHY4syVrMZAccdrXRHxgtTHtBWlFAM5iWq2+P357SLa7mDMSgvb3nXJlpUiZo1kB
VZD7sYsM0hXIPRQrc7SMqQ/Sqy+Jb+DuR7KOdVwQDht1ZsYAq5FjBuVvu7s4PLT0SfjjTGd8g5lX
H3BHNdy1vf51itRCKuCGqAT8wss1TgAoIPqrjLLQ4Uej+Rn3hp7afvp/Gjo+CHnsB6hvxeFkV6UW
fBO7moBa2agWUOL19FTnCXUBRrtVunlmCEkzKmJzt0lxr7vOXvVBfuL6Igg52gBENWKO0cgOANgD
gHB0s7+0pPMfUZ8rnmZe8sJRXmnr8aBHcEyhduFQZAnhCqAz5j3OJ7/YDNKRFh8J/wkCZCnZQqv6
lWV3waBd1H4UWXoLTWg1OPY6DyG+JJy4OarTWS0YE6hQ4l4ctJSY87tMoGVjE9Rj7yNM5KhQE4Gc
EIwF5IQD7sh8V886wSh1kOVUHdO63jQBqXozmyHN2RExNtZFCOHRMKFlRFxMgDoolYdCairaNUsE
G1wdBKBtg4egXpzrYAyVDU9EqOslkIJoTeqUGgC5qWBWeSmjWNGqr6q3/OJZXvOmQg2v1ULuBG+s
b9zzIIlsy3XrHxZZ51NWUPDHGXH3w5jLLIpuyVCepcjyHrajuburL5OvIg//O/RXPImTyCArHA3F
DWdNSBxrmqn4k05lbKGzSfaFssZ1LuMcmzuj2ftDeCdAtaT82fgb0S01Spfdn9DM1K1UBlDnoEiw
zgzBhdv0UwvST0EhdZxgIP1Ik3DQBpUDSqNBY4YIitXshxriiS8m8Czu9JRX0IK62d9X3D8vT3x0
frnjjtbDjlxS0pr+4JFA3cWPyzkJz8MFS+qpCZG9KEkiujm9aPppZRvuCnQI2NKVcPx3i1T2ZR4w
BlyDy5WjDf5U/3mp35XenVqKbimXQVNBJTVupZuFm4ejD6ZHeVfxFzihwYxzmX39MCyvAQo94+ph
NuSBR20LEndEqKqqP7lScBBPikzLq2WOFDn7P2wx7s2QK2ZiXuZiyDdrj2VvVxeRGNkQhPj6tayD
jR4ufKH2B15NQa2c0eSTxVnO2tmNz29ZmPwhttvkphLxsiQ92LT3F4bV0vPqLRw4ERYdxoNA2hTQ
JgnPMZnuCCsaVljR62VMZL54+WIZcH3v2n0AdUJ4XGTZ/pZ0X2dbCRAxzbJHWHn18UHd7PGD3lJq
IUzDvS1uXjc/A4mnRDH08LjLO15w4lLBOUXhkPcDtzfz4nE0sekz5uPOdtm3JbQMc3/eUDIjgv7d
Zt2ADu6SDfeRKvsDwfC0QO4xDMrYzjq41Wx6dB/lAITly2+uxMEnS8/mAwDR6CJrlrrJmL8P1kNC
GWwIuoUt7Rykk9jSWPb5AZ2nsm2rK4jQydLoqRWlWOloaIbJlYcvdVpHLYV4FTho0LAch8i1vXWw
c78hRZ8SkTvOx2FqAw3hr3n+Y9yFqQ5So2ahqG0LuWPB9jwH8lwRVopeWJ89WjppTtZbz8H/1jmC
AtARgRggy50BSqb0a2XGHaQ1bq3tIAJ3GOYdc+s+010mrxltkw90kXNtXX/iujRWJEfQPvsEW+Yv
OKQfB8QmDl4+WGvpMbVT5DdQWsLsxcNVhfD6t/WoybiO7YTZDlGU1hVnXzlw7ShC2hl+kkIxeK+n
oPSjGQB++KJNOh1FycCDrTSs+mO59T/ucPdwQWCwheCdOJjhFh7W4j9EEqGm7PWvoyMTrsoecCgm
Fpg6UEkgmYoXSKUCelTMKoT5Tvq1W83u9LS398FX5qWDeHYSnFttUtGr5ou7pW0uzWFE5gQmZM+B
ofJqhqJDVwxlIoBwOSmmgB6w+GqmjcTPBYqbB3DXkOqafDLp+718TuF80//nLUstWTwoHe+UXmb5
NWRRlio/cyJ87fGLY/9b6fIo1L2kFMum+8UbcCBYxSZhiiYhlpX9Tw+o8p6dbGDTgaohtz8Ew8Oj
TJSUj+1dLmaRMFTMC0xZy/wEfJpqPYRIDQaC1oePHfxbepJLB3UCrYZcxlHUhMW1ozk151XViYQ2
b17rZkyjpOFfANy/uYZ0MNIrB6d5laCw4bvmlsyxF00KpO5VjSTKjzG1yRBIUxzUDFML0pbz4mqi
4+Fx5QJpT1dFimKlr514VWeyl9cPyK5CH4ge+uIljGBNiDSpEKYfEjOSk35w/pjTo6jMQuxAupYD
w+M1lEc+2VEe1htWmrLdszHoXyxK7v3qxcHjEvrmBsh+g0MuO28fzx0StvcTpmO4Gey5IYFgwG7D
yeK0UlRCLY87UnkgoFp6VWyRFI3/KPpya39JhP992KrHsDPiTTxBagIthsduON0JztBSASP7vycH
2sq1q7G9yLjuydRlE06DcbRcCMk0TMymD9z3da7EKvhJ7cepORSYB8KZ5eVVIMJKRQeQhJ+m+6zz
lqBRbdbGTPGRG/zsaPOc3AR/z8PXjETYtFl3o4C3T1VEfjaEP2mkF3ZOcv346AOclb/jGsZX0yDs
tSxVHxKLfh1bTRib3EG32pStiGqkM3OwOJCdozZOz408Q/ZKj1OHRKQzbbffF0uz4DFvZI8fsBIi
VFpZqJ0Gwn8DOPXWAuWStx5tnVygnlTuEYVIxK/ZtTCswibS8Qvg0NfOOPWhyOtuNR8JX2FRn8E5
a9Lau1DFebVwaY6P/K3S+i2VApWQsZOzRIFctxTVeWMbQuRZhZ7uAG9JvtPDy/6tVzvC8NSoUXy8
8Oag3oPb0GDzdlCqXebXqUe3+R68cFR1pGG7QOKHhp6BCE9R6pYiN+NnCvnA64K9+64BeWYUgNbl
6sT7jHsowDG2BED7+annqjaIICWG9mKuCZEaAhVcmeV64yDE63FzZGi03ka2F+UnmtgtEKz0nuzY
jjF6oKziO7dNPuEwrGviJLJNR+ozOuoA/QhxqJZ/vrp/YlpHSXUKy1BMyrGWbbe0/m0saB8elysH
SnYMXeHwDyVQJ+7erojntYcOALNhOmoRcLnVgeP9DEzBuAIn/PDCTTuDyJH9v1DFZ8XHHtiP5rZ5
nKuJJggLv+Ni/hzrSyIa0c8EmgLzx3jvD0WjUWODg/iAkKpZIIzWGDo8xsilrYZqEmQ8gamfDVto
OwpHpEv2kOxJv8F5JXO8fZXn4MqlDR5vMD43f3wIYpH9zP0hlEp4GHYPwSQQtqN8nN65pxOogmeu
CK7Fu9WdLTxjKTyCNw+e8F9Qynq93tEFVXrau60C1ALCrgsr6x+4/Goqbfe2XT+MCNnnbvQF3nK8
vGQQmR9r/aJcU0i17pb9k63eQMvFn3oIbJtL8xA+cQQqD757T9OnBM5TYAp/x3JUt3oSSdEwAvB0
+vP3BwEcxlpJB6V1zCw/7LChnLrefcZ/IIVKsfdvwkE9G47QsO62TePuEF613ECugW1PfIKidqs8
jQut0EFHf3ntWoEr9RQKvGdzZ/I3JfhFMXaCHSKx/pJ61sXfePe4q910dHL15j/3ACzux/fOul0Z
M+lmP8uMSzjU2Y/ISidO5l/MdTZeBKTueaQPd82RZfRF5oGLJESyVP4TymMp1eTQ+8HHv0imeoOj
QI/9kUbMAeWLFPZTwLm9DyqPl479NVNyv6qgkIOU6QbzjT0vJG5kaJGtpKTriQIpKtMq6IsTKg+R
7tGzrFB7LAPQ9F5PAOaLTopYACmoNEv23a9HrX1UUnGEDBfHNrSHxy/AE6dV61tOStewxRnA+mwX
KxNRh4OBUr+ofJgiNY6e9m1rCBdp6wsAfiCI3Rk6Q62f3YL5B77sqezauSyQ/7uah5Q/19guuuUL
wSMyAtS7Cx5aggW86nQ3WK2GMjftDddvhjpnbJ8K91yvKF7+mIK/LiRCIvTLMKL4+W/qf39mTuoj
Quhp3QRX0fRMQSU9lI6Uo5gklvAchDnImJRNBsmWoJkuVXy/GltfOo7QPouA4nTfDzLiszmVwjSx
lV+J73YoFwCDKdF47ntbbGAX1lr04u8gWhoq3PRJCDCYXqaaKNpb2E3MLwJxd/82GcD+gblyAvyM
Q6IuQuA6u/ahv5wdNbmv53jRmSIAZohk1OCEOsh9WfGiXGOKJq+5U8mZ6SH5V9jqcvr1PCH1eKqn
AsfTEq1X8Gp/4Htgqt+6VBqJK5FQhrCauAO2ohOXqrNVj+/rs89QAz5GX9NRaaZXJdAaI6YL9lvB
/8gDDsCIHkwabGb1fQV2JZ5BD/C23W7At498Gc3Xe/JGSdgazcDbaiWJV1lNbmAs/0A/mzKSiMCD
K06+ugvnT1IQj9RN18uQc5fKqaQmarD1Rq2VqJTZyDnvsdKvQ1E9yLgK73dpWeCccWQ74ZLx+sV4
kupWjrsOM+tbDmkfwxLWXO02dr6wJvYqX0R0mrj0kVsDkc3qQCRDM6T1hx2EwBD2kR5HOU6wrnJz
HaahEv3qFsoE6nRgdyLRo5lvMognWJROpih60FfJenLZtMSSG8kwIyvfvQyPGoneebhJrMy4W4Fh
JBUFnGA9L0fmbuOssf/jo3cDTdE6N+3l1u0HHjaaGO0mjH1j9mNi7/ikZSwdgtb5oHWgHCIEfy7w
j+L+DZFxjEnJw9m1u+RmIJ8mMlhWqlIvi5B35DJ7p4bX7AiSTitni/t+JpFLB1FCzsXlqJxY7V3i
erU9h9H+XbIm+J2mZMukra2MNCGZJjenlOW3iUXLWMW79P6qlyBQ58zq7xJJjjqbEHXj7HETcsQX
p0SEgzZ2GMk92oqfCfnCTyMG9Hc4qhbpxKf77CqX8AjLfMQ828duab8j2aN188380NmhHVbwafIh
wBdUADK+DZ2QD77IsZC7lu5ffmalwMu1DoLj1q9pCA1flf/wXJEA05yMH/nRJjLNxCMP2Ltf8L+S
zVqvjb/pCbtAijUx4uovBKvCXfft5rUMEgDrJOC2LH/qHbQte1F0f7FOGw+d/45dVIsNVHihIEOD
VdW2jzOKeevc86wprX/o5urW1gcXk9YnaMp3BhKdkbyD9bS9fWYlnS/1BEk8YJwTLWpkMS9X21Br
dAxx7e3MchzU1pzKbhPDKmc5lGHoL3v0bZpzMKGaCMHSZwOLaOfvjLv6R/uIfNcXmDhyhOJtev6K
+pQdjp7ufIRRhsRGow/DiWtQrrdMJXrX9l1ErglbUyIxr+JA4P9MD+/UvGTq6i88FV1syxM5z6gc
tiACeORkG5SkSbvXA77pPQsgFhtZ7eWxKv8acf4WYuoRyQ1++COUyq5cCK9AqCLAFueavsq7Ltg9
cdtk+TILQfAbkvbI5s1bLHilyYiRhkyer3z/uIHTd4phHTQBhz9hYVU2Wtq9v7HoiS8iYQJj1DyS
yUzaqHITfbEU+uH0Jc4OHU6kC8xpQL3Y443mHHyPeNf+C3ddVbbg1PChL41LheXMePWYaM+i/9/G
SUQsF+BTkHgohBgxvujKbrq2NkPXUICHEISGQtXDNbSDY+j31bISfnHqp+z6LgydW4Wolej1iSeH
85edJlqxSegbN27S3EGUCChSL020T3c4CHCOjokHOo8yuVgFrYABj2fxbHiHsJuwvj9GaLJklhA+
/1gu6kADWbsHht3aOHB359j285eKo+bDRFdqq9eg7RO3lZ+GGBP8lLBHssRw2+66OymaIYhfsCaR
ksI8ZumceVhy3Mf9A2PH6FuMxDzHh7aSGRYPW0uvjxF3PyuNOXFnsldGfG2KggrmNUqSAo1iCMbO
SWoO0TYp6mUoc6joJwOLCgUDpcdebZGXnXf5O+hyP/AYxhzoJVZgzul5mMwoY+k+Kk0zMynnDFwp
QygFnGW8EyE3XrFLIg2MeEQ9Lo+6L8coF9CavKwH9EOeQP8GTZFDUwKjnvPyiDlULCyiYQt3WA5c
fjQTrzG5DLvnDeM28KXhkYj0FZmyKZ+8nPI+7lX2s6YuuyQUQEYO0x4vF+w+COBS0rraBaEfEdlk
w0LkmKsP6PR9qWyScn4TgtxYQHnf5GmMCNxjkqQdhSCmjMJs+K53CEXe2old9CO421aCBlYMO1m3
RcuHIYXlP/Z6vk72V+fRry2+iGipocgq+eqsoeJzXl1mPs8+SQcP1FLecafGXOUgZmvXlqan2HC/
Q5NUmL0FU6yJZuP03CTfLRg1dZnp9evGVkDA8Pi2snieqWkUvDf2h4KEFler8dW8o8if/YJYLNF4
hTigVhVqG3PbToeW2TMmixrM5Oarss3XRclNGxDM8GY04cN6nQj1sDM2YaWdwK/u9zhJ58At+Iz8
OseeN4tCXoQg47zznjhTUI7lhTqNXuXoiP3xnuntxdRW/uFkYHvKZNBEStRCpzLsbIwv11WoaC/P
KpxNH2JMr2wMVrk9DZrow8ObeEixuN/b2wQLFfPu0b2cRTNEjW9+2JW3E2F/3XRl3EjqnYWVnXVU
TV00nnILDxcl9RfWVss/eIuWL4oTFIYN+/jr0nUTwHXmN4WqZy301rIvCXrAZmSwqwis8z/X/Uwo
3lMCKiOtxYEXYrqBXpOVVu+SNc3gUoil70VlQFwfcwZBRd8S2e2RFAEbf7ZYPNfCFglkHB0KQ2T6
kkynL4KKSJ3BmMCL/RY+FdFbPtKavBvGZQxMnnHl7VyzrHjgBG67QZ9hiuXLuBYXNqWztseXOe7O
IR/QKxsxVmPxfNoxZo1iTXv2DHu6Rt6nrOmNnn97+1ZQeVpcaAU0I0z6AL5kX9UjShKwOjmyGmHO
BhJpdZynokFsU0xwePwLsWPJPo0uQMFGewLhNjaI+5UYc1a+FhEt771S5Ji0W2ZaqSBJfr5lo+lN
VUqrQb1p31FM/3fmQOCSvl87NalHq31IJjGRwkR/TNRYHmDeMT+1hFt3iLAJAvT+uvLvycCHa7oK
lFr+tOPJ6jr0wZjM6pulv69HGlZXWPMIlFDe55uFx6ptNVInY30kULe4pTAkIhEjntNJC6HkCpu7
fDKR0yfhYFziEMkYx4MoxB9yOHenx1uX8rAPe8dZFY3lkrE3eATVCR6w66G5a2TAIkenA4KuLyy4
3VfTgUDkNvo6mFVG0sqHq6kpiLbeC/gGayQa9YlCNwaZrQhoBh/ULSfXZD4f80lKqzG61m6N523f
eH+RDCvZzKCbQWSD4+FN7RKlTt79RszlxB17tk/lJQbR/r0IYEn//XJ4TmMgUpEGOPDl7jOBYAB3
BwFih13w7IN8g64kqjYLqvlMIQkDv1NIhpz7bvucKXdhTg+BA4qUqNpjrEjngzhdpFclANclykEy
U8/sd8Zk1tOBf12Uav/cMGe2xbXJNjuHdcQztALQvKmGmXZaavoGcefw/QFY5hBTp3WuzQOVMJpd
ZQxV1iHYYGFjOaaBQ8m7HFJ8qGGbfUILb7DWXhxQDhGy1ryc+79zVRv8AshS35H7hNQRanmMXh9E
2YB6L1ywl/QrJbtDlvRi+S2x68p8Nu+Lg6gbIipkG/DaeyR36dxwqBOjZASgjOiifbww3fVCxnhK
VVqybLhtSN0+pycOYsyM1WsddHstfXxX3qYwT7+4v2OuT8/KIeS4J6zlsYL+E66zJ6LelAUQRdSd
wufvLVoaN57RqNnsQAdwfHkL1NHieofPtuHD25oHgY3h7oVa8bBFmLwysYe2gj4yF/aMMXOxJfOa
mnA/xwd8G2t2yxvBd1Mx8SUvo55Zhszbt1Ghx2Dhh0es8IPB42KrkaXkziahYY8Kc0zvT1pG6lov
CydsWBI0elJw0AQ4AlfM4LNhIwUITumvrmO1YFW7JkZXq9FuM2Gvek8gFBhTxFQisNNpS3f7m6UX
uacuLBMXHI9Un3XeYHMaXfStQfEo3If3S7wT9wMKOyxfs9gWRQVSzlvRGqYU+RnyhnG18YpGSObM
sjXiRIYBFdRITwbIp9GPqsdl9ayZKFmwsji6iE4Ve2vuTuvA1kfKPmw5QXNeeFXwmqQs9nCltEjw
8CGqpgdlv1Hp6Cs/J2W4mw4aPxEwierz78MAzvDVartLOWaTvpqVYrFMt1Ghy4OkOXabK9AHbi6I
dQ9AuAQnnPX98A73pcT64KD3Vcq8pxER5uhUBbKfSmOG6hJq0iPkk/645DOkWSpLm6HzKhoqK4bB
PsrGjeNCTLsBbGnfTafdhNZO7NAbo3TsJxcygkk90aXgVDqzFLMkI8rMkpXF2ZuoEJ+R9wx11hfb
Qo5552kri0z0meCCEiFu58uUkkzGCkz+lpnt8WVLMOuEXGBv7KiRF18Jueq45asCSYVlCrbT0AiZ
zWmBmhA+O7IO5i3Dw3qL/qs7EV51wpWHFZPGBB9AMsccfqhceoxN7vC7YgfY5FNkW2tHCRhybZGn
toC1Ez6oiJuXdy3IhZD1/Egfliow8CjxSsxS4uIQ2a/27u+Q9+cy2wPSvFtpqmMDlX+XNFb82Q5d
3KpDZKw78IV1N45eKpH5cRsyRUEqFUBW5F8xIYK9KeVzSx5Nap7MosK8BTULJf8UPTn6Ehs6OKmp
q0CemF41w/UYwmQllRgpIHb0Ckka5CfZRz1ol3OyjlzxYHeupE2yMOAzXT6W55Gd1ObOQGfGEyHQ
NZYEY6xrDYvcoJa5Leq3guroJ5Iak/C2K+Wp0+0mel8hbujXbNRVYKwIc6MfCIKl59NZ870kqgLI
sxcUdSKZ9wb1erTC/0xVLn/VCy2dsy2iGFPeH8T1TIKKSBGFNMUX9PbI00RurQf0w+WQoi2YeGVH
FfaXtKQDJvBS6hU6h4Cip0fXzC0TAmRjDUXOwJs0sGbQfohAnQekr3Iw7YsKyGC44VVz5LBlmwe4
g+M7DiyB+R1pTwTNRuzIzd30/1jc2IuaxRHtNA9n/N4N/ra5wte/7hFzX6G9Fo99x2mWKSG5jrn3
bSbxfAuttvBPJDXp/Assq32TMESRPhbNnnT2PNalflPJA7KsYAR7hZ71GhIJg0x2yoNceAUxzU/K
JXt6cQh71RdCOIzc4zY+DnFKmCxSVWzXkqE146VBgAxy95rzKtCmUhm73njliS6yK3F1EiDGlLig
LHlXnQIrWb4ZmHmrCzKNXn/N0iZ9oOtjNG7sQcISObHmFSdfzDl2XQFp/ZPOlICHnC+/0Lim+0bE
/hjj8469qx/yxjJC9Tw7u4YHoVFbKX5GdZ5RDXSV7YcgCcsuppXo6xt08rfROI8SQIK8Xazx+hdr
L+E0mLJ33i9FwMsJ4yHBznMkKCWr/Dykne+5HDbJYfC3t2yBw8TQOEOiauRmzU2vIcpQF65XLDsi
ic4URkaisWj/xKsNGnhetPlbUQIUFLV+obcnxQdK1s7qp8yJK7RW1+oiVTZLOCpIGnZ0e8ayImkK
zuexdfGM9DcOhwoetlHapAEmzDhFNHDPlNyfQSVQXxVXxGTq+FtqOO1AFYDct0J6LkzQ9YZXGHH6
fylEIy9NADbBxDQ6aPCfPBWd0TxdXi7FI+AfEwvNvN62/zCjF+MsP9Tmto644sI84Zh9miG+DBMO
MlOp9s4cqfNII8XLSG0Hiq7wSlfK1lrPidT8DjZ3VF6ua1WErx83sE1FK5hnmod4fgVOdFTpRvqV
Bv+m8b5qpTFSl7AGsLfRTjGqRQIrSSFB3A2GgAM7TiSph4RZxylI39fG7T4rUZD5SwZQrlJMMay2
8NEQdNDdF2tLbCo28PVSiNQaHh+T8ztp+ya5XvSB2fupPsg3XKKkWEsWAfq9ZCSvBF7hM+IuwEU2
kM3bOg4/m9akIg6yTDffrf5z+LwTKul5p6SDvTyHKYWx93Ln6fuT9x5a3xgwqWOXMCBWziukvruj
wVnTqAdtX/0nnG+p//mKu8YBq42ZKKAGPk551juAk38Wn0THFjfvZGP19IRk0cdjsXmzuIb3wDJw
DLF8dfYBq3niDNGNfmGNSkaxwL/I2njqobPb8sWQc2CA1VGgr2hPYqFeKjv+8r8u1XcBlR9tX8ex
ivrO0H2fyuL58WBOAr8bG/rH0/XUbNsdYgIt3zkXHN10yyYJNdRNqz9Nm4xMYPcd8qG9t0yhO9nl
njKzG76ekiGcXiNMjDPK/hqF/kjY+/hSbrJQZ/GO9QqsCsmxCeUtHCGcGqzqwmaRHM+bWU8KL5Fj
rtPmDvo9wrsRsqx66FjfYPKxGWVEgr6vOq/vCcmyxe+iF+XycP+LjhsTpDzjLyyIV+27qQ1eeK43
P9joovv7yHt5XFIx06JJ0rQLF5Q0X9UhFIkDXupeRP3eWYHpeAyceKDDZtsq8xfRpCHzDrkA0GHT
qZT3k2wq8BPISr2mA7HiH+K2j8aZ5Pi8ijML7/FkXPsgdxwRc/2VieQGnA+K1gge8hN+Cvtfzck6
Mh6fZiUn6LM8VLy3GCXc8C255wD6CCMFDmUNRsmknol8AxT72GqC3MsouuG9xxGhtYeVkCsA8W1c
5s35ONb8Ov4QNQf/TY/RR9Gfm2P+1FG4gE6azZaui5A3Pwj+N3eqc13PRlL3gD6NoMHhbTcs/+LS
HjkB9CKdHlS//iJdwxfHDqWg3Nj5TeS2ig8h8P60Eih9v6GCHLwq8XEf50VNe6uhrUDiLFbweFSQ
LYGrG7Z1dlYRMOflhzmuMJX0hi+5G9RlhRGJfqTC0y0O7N8F5Rx5Tp6tkjsX5UYNLUFQF0eUyErs
01+SQEYDEklJZiIgD1BE3Cnuhe4rt9/FWyuUqyX/kPMWMgbCySu1m/5Q1oBNtH8cJ1RKZS8pd4t8
BCmdRELr2hbELO9tLMUkm6ag1jK+of/6s2Az42dx37eD73yiNtfKEtQOyBrWgVQouPoSd3XtwVF8
Xa1uvv0D84LYlkAKIRLoW5LJIumQZ1Tr9unr+3s9rHk8KXLbJwmxxtpBiw1WSk9w7SmcOrLT4zg9
gOJxblauSbfuqd0MT993oo93k1BjSjgIU4fTA3MvLxOEoTCub+at6hVsLlwrXLxJH1XLt2tX85Zw
a6EveNg5QXfklWaS4n0IuDLPtQxZDfbKoqNsIOqLcPNUew4g7BhG2Z8ZPzTTFNy/PEZafJ6gylTX
xX7mm/nv47M+CEbwXMfRL5PiT+SkOlJzxSU9pYKBjDcZNJk81r2DFi//z9RKUHziLcfN1/LNMVEu
/UnbhXaCO/sLDPMUqB1whkNoSA28s37TLWgIgg/7h4YfRkUne46ue1JBZE4umBKbsw0OkQ4KJcIE
+ZmKBf9emVupAYod+y7nGCX7YVllB9DfWcU9bnnZMeHLTmDF55bed5ndz+Fx9iMQMX6f1T0EBSko
3R//gTOWPvmTwtkXx4WL/B+PS3vfGLLyN+HIMo4IDCPBq8P+KoNpuJuDgXDWSDhebVYXpD/sFJ3B
nGIBBjj3MD/QQd1m//pamPklOZdR+QdctfGioZ56AhK2NbQ5sKTNsDtQkk0/Yh9bMJYL3u6hPH0A
UVlgUOEbCAn94rvq6nzU+ayeWWLBDqXgMBhQuVipx9pJX0LMU7ywIoTAHJc5KwDesT77YWImhy3/
99CuR/8pkYlLdjTcXeAn+Pm8SBPfmqTEONtiXlkRxNNLHD52Q+kBW7catITUf/ygW4YzhmcBk0kD
tCB5um+BcvZ5Z/e3nhYFSr1VtUDfJUXgY/3EpI1PVGiYtkveHUoqPdr69HFGyBpZGzHT/bhnAiRD
5rFbCEcqF5bRyO1x+UHkw+hnAET0xqzv1GxG4DVkFkbc4zZUBm7kf8BG1eVxbwds0l6RxblJzPcY
a9ZK3tB7vBolhZ25a0uyJfl/EnfAbpanW/B6jbV1zgpbXG4yHr15qfUi24JaVNmUtlNW6d5ZfrYq
S/WZhQv0P2gRbLcI1/LJReO5gp6m/wGZ8MatIIej7a9xTH4YzzSdFzaQ9e6jE/8KINIHBc1PUwzp
Wg7qOVxeD5AT/PsCtBRmK33zQ+lNUXyZzNl/NJGQ5abPhoQOCti5oxSRPkJn7KlTQpnumEJKjlg4
EZyOsOk2Q8AE5Pzs0vwcOJ7ZnZKQMkHTO6Ihjg/wIwKjuvPzU3R6Zp1bCZ6694npbvrSI2Od75jD
42snAJEkgMgFsR+YYn5sRkJ3i+oa7WTwlcNLha4HyfJtJIkUgNF82AMDKlKz6SfTExnHYwxZtyvQ
F9HPwATOvpBzRcBL7G02RytPuyaVc94MNrs3WMf6Zo+SkydXs6PGmzVytimIsabam+UqQ1if2HkY
DZCIwaKVl68ZQ3R6z7FVY4TbOW3anLn/g7FNrJiAFb3AdC4r756K27+utd3VPCNFYFOGpY7XOZVo
VlDegdNf71ySYo8kVcSG7/YtpDEfVARznkSmGDpKoEODVOxYihTxKAS+YTf8cOGqbLtNXzt2rLsW
mBik9IvjQ6DpenpA4svrffbiayRTC70/7vWm3qBdooDF9Fc4JLJBTyxznlo/rYZlmE9qKF8URmwD
BXzbrTuKTFzZy1VhMKB7LeOrlVyy9KUm+jq2RIvW3uNsheJAJB5tnDu3cTNGCvSy0/9yh0MN8Dq2
m+RQJNyJw7wGC5mkdNasvZGjLEgrg+U4rgagBseOttgqC+EXEVDnT/SzQOB7oHUOd71R2QE+WCUX
N1Ga+WYSP4WxkPwlof734Rv4TSphNSB/s4w7+tUBYf6lfvV05n1g+AJ8qM34QsPAi+vjOycfjzdD
il3TbFenxVygBybYrhmtB6M+qNpg4LaC04MQDC+DZowBRnJFU8W7egbp9mDAgXMPjCuFaHXXg1Ml
9sINXIwq6JSmTQWNV0S9nfoel2Qbh42MuaucD52xTmE37z2hCzy7HTGJjF/xU8Ii+2x5M+GWPFAW
tqqMc+oJXZuDCp+bXjPvzYaaR+ONlk58iomDQUMAIED8clXgcLXCfR3Qy1AVDIEf0PAaCHlz1vov
E5ZndmptkPFRhBkMZ2jyQYEa7/4jKjirrbPAWLKjCyK4UWBZhlGqGD2Fj40HK7wna3jBADiwk3uk
kjXDKDbtqlj7TeZQM1r09f8cUG5ASSNVhxLIVaJJTXZytNhq5F1TeDMLRg5kUr218cSZYFHIg4xT
Nw3HigBn/iQW+sp0Cqh2LvlE9UuIHZym2wQ8MgaE3LPiyyvO+uyqFAeL6dqT2DbPxYuOrdOSDl9D
UP6Lt1JVggYzuVVGILvrVwCoH21xcSEB5GF+YkHE6TvsgA7riAx1tL1eA1AyB00k64AoGo8vjS+3
kajPFWg2yhLwJfycpG6m7oYM2hrQr6UlaHoci5NL0O9VGLPLUqYPBx4mkEsFG1sfUGKgr82L65r1
HF8HMO9kBAR5GGgPrzv8673K46hv/c5YWsEODxPONad1QRHIa8LWLC03Lp6L2yDE6FnuWgqN6s2j
eehl04XMvbueymxDYdVVeR2Ig0pMay44sKQE+f16HoDeEo34IL0KZBv/e30vdcHYo0VSpvHA1Htx
zTOBfAiNVUl13lFgND6DzPcV/DCmejXzsLMfEHdmXL19YbX3FKbrtgrJ3z3JEv2zRdsK3SAolk26
tTP3UekBD/P076P0XGfFFhGbk9yd2ouLTKASDAX2cMpCXsCxDfVHwCGNoxo1QzAY9H9nntrgo3va
0vUQozVA9aEgfslmhFVU4Nq8Q8yh57j2Zy+m/glzES8j1HE5PF0d3a57BhV5a9L5g2MCkb+5aCW3
sgz+VP2RmaD7yowysKRZFtilwmQATQ2NrayZIeDgEmPK6rcXiEtWd+Ke4+Lxe83uMMXmHnzMejWK
rnkKgxgS2j2sHEndny1fv4BE7FMYHy9IYIX4jE2F6vm9WYri37rCKbKA65PoAD1wZLLtact1LbeV
ugGBRUj3VGEoDPT1as8sz5g7DY0vZx+izB0kTr9BTdtlNRY9IpBEPDmHjmJTdIFkxXa0KgTsrUVA
d7DfusGi/dIX4iVcpdvfXPnbpLse11VTS96RJsxPIzVEIHGrzRXOh0IuDgtWESkIFH9/L0cat0OT
ypRFaGVEFMkT0N2nDDDaL2ecfqgV+UduJbuzYjkWq22Sr3P2VFyw2ODTAXXaGeAjqUnJuhnvDqdD
qV2HIU4gzLJlp0XCTqRydupoZGnqj1ZDU42Fy71UPbL+ljdgq9VmKuQIuPbxlgBZdPULaagm5rcp
3+RrIQoncGoRLSbJAxOh4x8C48hiGLsSXD78JuKLvx7OfsUHqDZZeNHzCv4jpWSAxlTWh0BttbIO
LszQ1gYEy8Xm5J/odncdgofdteB5bpwOakzk/LPjM6n9Vsj5JUl9zduuFFS7XzO7efymM3ZWehn2
HtFBnKGyPqKowyUnjuu+WGEV5ay6ktVsF2O7wG3IrHkAy77pNRLDNKu36TYZ6akv7ZFXp76z1o9j
Hzl8AXRjQmuD2V1aUt4/y3Gj3xz58iXN+8+/ylCH2QmUonGXRlElslxjjttdqYjabdX+P5nLkzPM
gAhdMGdkX3Y1GmmQ7Rtpm2MLvxROyD3hP1Q2tR5Nb04dJgKZ4q6b1GlGFpxjrsun+pvbo7sFDtUT
EH/oyONg1BnBCVTY3VSxTh8xvN6pga+lug1ESn3xuS2Pj3frNETbMVaW4CzsaQfIJNKGA1bgN+zp
5NjiD9fW+I+PmcX7MmwHCZ0V7lwiemMDy9T5e82RRzbDuAuMLk5W+Kn0iKNJlAIAoe2BD9QZAuu5
BcJxItgCDwICN6BdmePnz8rUP7Fvaqo4RSGtb2X6WWgZSlcENnAFSK+LPBefM/Ql4cyikW+r9Dcj
por7oLVsYJYZbwmkaWEYcL75o6jQOx3ZNY1bwA00gREME8EK6KEhXJg7dt0g9nO4Y9FDqag5paj8
HiIxaBXdO5Jiws/A0nsBCq6S9X77w93JQPsVrRwgT4NcnU8t5K45YygRToqwy8tNrbRlcQvN3H8Y
ip5Sfa1uOkODK3ZD9+CzSsHz7/2aIopmvudJagBmWUvlVZf5OjzgNMPN0s+whAwkvDZRKB0B1zE0
wLAnBqU5r9v4f4FvlnZmE4g98PEHmuAl93D9A3oeZ5aaww5V397v/xyGcNJDVGLnd/SCX3tWIxFb
UEaRpGB4wB90rd0whVS2q9pNs7DieTl581BHdXQN0nmMMNbEzMOZ9NJZx19GDKLXeQKFPGOMWrDp
bXslK1TLN9rrAKxF2c9kCPbva9OsEh4+CPR6k4jPZ10ySHXI+pZkAWvU0K/4nneHMlFX5+ao1vV1
tiv6exxd/DwOLgEdE7w3p/gdF9b9ws5gqszgyDjpg8DGCpDcGLhu4OmVR09gg3WBZOQ8oHZezSP0
tTH5H+xtfehRD+o77Zibc99B5GV3SuO0l5OdnxHAgAOGkmaDvuZ9MrAQJwFvLjGaQ6Kb+fvMt/V9
rKtdQVNHka2h+bOixCNCb6//kc4Xoh/USzAVHGfe3T0wz5uU70ziiiryuTaody6vLgP9Lxlgamp0
vQRzLKPkLIMwQ46RrIZ1eMIu4ljUp4L2G1uSKMY08Qn5H0+jGYrRaUtV0jdOK//ky3gRghtQXv4b
mdL92bga8udVmJBZIwiQFV0CB8bZc5abqPbEy8MFRR16jEeCREqh9RFvK5sBhTO7Z/BpTViLc34Z
mdtuMpueKgcWRyKUAqeY363Q/k00zTb06C8mO6pp78Pf+XDS4N0KIrVXt+skTkucEKTujCXZz5cS
IwQ+K9XOoSVQyyKcKOv0+5nuxzxVmv90PAH7fhYHk2TpT8g1PELHhLkQvDuRfbplar2PWPQ4BWBC
5cViQQ3QTfbDiDM2CNOWqTBvpNU7l3ExSU7hnGDQPOWD1CH2ADup5Z1N8J98F4y7Fgnx3nJB+QK3
47vxDES/AdoIaSeovMADyDSDz26uECTG1EwOcYJzThzgqEzMqENR7SyXqnUKzTRppz+kHiMSlCFf
xewYpEN3olyaFJZIIo7GOCLlO6DbtRE1/7s8WWWQq0A1KPHN06MvG+TkeSxv9+fy9bKYSP+0heP/
2ND9JdLz9W+4OnbjV+BeEAzeg5tSqavBiE2mfZ6Vg3VuqDsPGD33r5SuhN5TRcKw8GdDYXT46nyH
EgyWFbFhnKfVXnP5RmxLvYZMNfH35cENECOjIERaa6VrxBWaUFXMPwQiKqqXfEI/1J+7PjUu/YKB
NwqXpkAsRKb8w0hD5422mLfgK9F7IS0xTxJZKOUFfUjx8jpbIDPnzVQ9+YQHsVQG+yalDSiEFaRg
TVsqpCNFRkhSyQi9y2/0GNCwHKfSNDG9ykfZk7GmltpA9S6kGKPxsKhOGcMUmfxF77r/mnm5MQbX
In8tBUONKX4oVA0wV9OlX7vlcFRad+waKC63FMXqzALbaVxIg6zWHTclF3kOhG1MXlTeunB3jYgA
HUMGkEubWmnPoO7K4h076LzM438/bdB2airg1JVob26iMA0Bfplr6q+XjeQ73mp3+KrUg4xzuNys
QvvXXzOpVwdbqu1u5zKHPWugWkJp1kB2Wtn81mmy/yoTqaJAySK0vwb7qSVFpr2u8FVqF4eTaxQX
mWPNLPfAW7w2lsPB7zR8SaDE+G6mNYTr3zjSsSPOF2HHRP6CezEUCKV4m9nIJoDxnepKSc23YCuH
uQcFmxPr99Qez1PM8wPDvebH46mEypqAuv+PO1rDf88Nwn/wNGMqerAg8tduHTFj9Ble0s7Huakl
/w5fZWtG1HvLZIPAhHye/sOlK9AxqiK0nxzHcrKq50LEWFB+UquUElhlRPi8tJ2OqqVSrvjhFxXf
psCJkVi+aTc44JQei0Pit7IPS8jLmmiKvBMAkuSiHehNaIad2gEXZKRClae6pi3QKoGLCfz1rxDT
OEbz19MKMnIs4Yw3DhVvvUBuzQERmbSVwXj+1C4UnA8sEN/OhJIVhixoslGQUUFtqePT7Blq/wQv
wCQT4lq62XYKds1mU6S6utxzAeTexF0wO3LVCvGh06y82PmPKg7xqN8mJd4lD25EzHghHSJhkOvB
Xl8n3hvqKqqbP1ztG317lMovxKwQqvr/u7xXdL2k3VDyYeHLzwGk/Y+HwjTieQBwlvTagG3ArBc9
9yy5txTM5WWQkMluZdVRwFR1g2UH1Yr60/3Gy+1XrsI0Oyr97GvUawCS+JnexZPKwLSI9IlLBt72
zbxXC0heUmlAfULXBTqhYxl2V7am383wnEutrjeH3E0E26oJSHSx9qUkmeZm9Vpdh/sy9ywhoTIG
+TstYuGu/TVgr1+H0wHVBZ651WyMPWARm8UaCKdKS7iy0X5IoEL1G4e9p550N4wcMY0NQm9lBwF0
kPjCTml3dpY/bLsiC69xC6/ibum0178spjIkOFVCbyFwKVzmP56f8xBlHPSgkoriqxV8EEtjdPq4
9KS1XgiErJmz3OUOb/G4Uh47t3tsW0mQzS6oEPQKSS4oWnkouArYmbvXBgP3+J3ik0HLqsMwS552
oXDNQOnmA6e26UmLIhI+5jk4KOTqdULMiT4YNjjPDY3oYgsB90OtB/viH60YTcofeD1MthmMCG1F
e5IAQKaMdELSHozOMph0NFOEmN20GwXewGzDn6+MYUPN4JeQJnpyLrdrmCMvuWlOnXkJIFmiv9zM
/GEA2IY42soin3Sv7GnLwG8O0j0jK+egIBVpjVZI9pK7MyefxdgYoTZjELjcwdA1A8s38bRPbmNA
A8HsG7WA//Z47x0zBzObKv+kwn9CCEFnjNKK4rKvKf9zpnw7jdgif4eXLrb11VMGLLLhJ3bIeW2F
Jgit3+79EgXv5HNBVfC97WQynBXi0zN3KJtLx5KJfoGIz32nkLQZC4oWO8HbjhgE5XUlurxn5GGO
/6MZ1d8FHPkJyfEc8rEiwz7p71d8P1ZOwzWAa66fFI592AVFATjEj302dGNXZUwr5NE6gPIHrFtp
9Hcau3MKoCxNDbtCIlUjzFl901zK2kvaSHzKaRDGZDkSlg4mxnZ+NG5qicA12GfI4afCUcZsVgZA
96RE/Qkfh8SeplXHJ+B2nRCW5jDdEuooVXxpAugPdlxIPwgGji2w4VxSOe3+fc37SlOoxwXGAhAM
EcDZgCUsGV0ShRiDzZC9/M/nMkGrNis0DsJ1cv6T4grhMa6snMpuc5p86hfEc0nXzBAQ3BcCWId2
GGd6v2aC2nlI5cGQBLT3Io2r0WJViyv5IGeo804IchEDBk4KDPted187WaMWneaSa2wbq76vZ/5V
Bv6ZBxGmn5L0W/VbAQT+R//qTkG2b/MFTJiR5ERrH5s47phBoKJrrd4Cb54zQV33YbzOWi6W6DDE
HiemIuLSmgDYxYtZFUrXptoIXHIMZHJCu57TFGM1/8CFrKCSJktL5vQiSdiQUwt0aPeVGXNz9uaL
tNRcy3dJTvHrubPemwiRU+9UMsS1Dv+BfAh6BhKIKBhRTJnNd2WVdFjedGx7kiDRtIRybJKrzL20
BFJCeDujfgY/GLxuwMZdRr1xD4tAO5AcGH1yQOSE50De2yqY2vuwP4SwP6oT/wySnQRR64TStgjd
4SPv+QD2WDCiENP0eYMDd+OW49vLwQYwWp/czt+CSV0YTLvx1Xcb9rp6f42um+50KftqpKKILOHX
S7mcKGUeQqOCUExUku4yQtq9pfgXrsnp7AMNak8g5QnpV/52H6HKG1imAqmss5MTHvQbFQ7dOsWt
basKaMp05x8f93kgmRDLM++4tzmVnCkXXswPeCGnSUUMkrfdc7F5gEqSU+4U0OYH6q3Ny2rFzf0s
q74ur9e+ujXIIa0m2nOxazfigYknJeBOx9ErYiXLaGCJgFr6lPyfDoW7XyUPtU5P1d7ORbQu3i6Q
BpJb6q3BeGJBi84GnazQJPygB6ggpub24tvTcC82gz087bbUwHfLx3hy9nVYNluq1nqFEAUFKPJE
qZHgemg2/fVW/4e2obDM6fXTM8k7KaPJB/cm0t7yOFSN7tHhwSmiRhYwrXSYiYhhT9jKITtOnYgD
XEQqxF9PBSllIeeK0VCnB99RaeXn6nd3aYYH3e3IuQhwsCvaQwFxEbuVJGCduY+79l9VN3lrRipj
28HnqggVQ76VWYfSp0WcAVBPG5/WGGZBlQq5+UpjIG7ooQyAM04R7mBPimh3u/KlWL0PppXX6m5C
7oXj1lq7BYZr9d2QxgeZU9PSe80l6xM2ZFxTuxGbcgfkaI7vtGWJ9x2//rUTlH6uDUK0Xjxsygku
vT/ERgijx/k+Y3YIY7/qGjPsjwJ/BRbeEwHGH8cHA7PyZwBWRtWXIMMdNpWqVTvWABySbfV/OmD+
xxDnNw4FYzr4k1hooRmZu4wcVTKkgVNAqvFttyhV3g79tZVemMCwtoMv9NYXpWnrMs6lazqvRION
tp530Alx+84ORUgHWBCn5nW50CJbT8nIEI2A+Cs4Kkr7s0ylMQ56h373iDLP6Is92VxTkGxcJOfd
JfxRue0GNLLnjysIR7If03SVdqjVLVSuWvNbINpR3SEsTKy/bfpHWzrt0HUmtZN3wt0GUCrVcsAQ
13eLfl6arpv7HlR3rRIkS0JIi5IKOgLdAcBDr86hABB5kQknkCjE7hznxRsdvBUjs4xp46MunWDk
0J0KCUFceXA0+QSTWqjMIkyPEm2G6pmhUPsz2I9ah0m0rovke9sQjpzeGqGzEhCjjNWsRX0ebuUd
7mj7Vgp9ndtyyY77jD71uxZ4+EbzYYE2ATu+W5ipYNj9Pv7XNJAbu4PYsaT7eDh+Uyr2Ke+5bseJ
SIIYRtNZShA3Iy8oUQaRGEu0tXXsEujS4Mx1K5mioXqlERZMi8JbTwm4PIQCF78kjzezjQUE8siv
QDpdY4VzFHrz19vmsC/VQSz+xj7o+bFhdVXu71Y1tzWznMZL3Si+5NQikbQYxHcVv02VRdp7Nt+x
wNu2fnql50N2u5CBL1iqUosVg76W1Ws0g+pBy0urpxUQnhmshPdFmBC0CG6w0BAqoWwq0HOSaC5N
ViJGSfwl6G4Q0mtdndyIIakku6y+Me6f5sMX6zBLXem7LHl3FVF4U/d9iHEtJ64Up8kxO4GVTYsX
llrevGx3fAyjP6G/STHjEYZi2OCWH3TkuKWCj1SsH0UNDVgBtotfoUf0C29hMVf+rLHpuO3gQPhi
1RhAFNvkFISDXBdUDSB1/L6TtsqahJg5+uu3lMDUU4PvIVLbnk1dGNhApH+bvYtCfV7Bysx1+s0a
k6j/4Ko/VerI+ZBRp3IWf0ZUMnEfTKS6uf70oG7/JqNZONDH5VSccNQw7Eff0NLRkKOduaJWV9K4
a+LCoxxXVcTkTUCrYznVk3J4oRjlZetFUwk/sp8yMEi0kkmDdvuPzDsIheBASE1N9QOwPtzfLoKT
vjdIwz5FQLQB86ZTFPiU+bj8eNDQgBZwwjn2dPViLv2JXRtjHMD6tzle8a78Vc8+ym2vq2l0B6fm
Ta3DcnBhb0udjcOoLnGVLeWQWgKBUpqAni/HN2Hu8g/CoKIYC9OyuJO0vYzMYYZXDlId7fJ2bYYz
OqRuelhPCX47z8/PP+MoomThjqS3e/CgWc0DSKx3zV9uD7m/c6UX7wWkOhd9vm+nDSjqZuT52XyJ
8iBH05wReM0Zz8Ay6EPkeeQG0/y+0wc+NgAIEv0zDuqwO2HwnFtkCFEgGVI+3nr5W10+2cNc4SxD
BamGNc/Oa9capJWOheNGEbiL4cjtJntF4pNyNhAxgbpNZeY1vm0ib/Lhl20WQ+T/rJFWapgLuTko
8tuI2HeeoayWz09SZgS6tXht9OEYqTU1Mtkdy6LCAhXnHcFzH1hCn4npy3NhxAIl/lWMj4iKBWmD
vrSbtrKpKjSdO5q5kdJBl8KLOHAKGOzGJ+7eST3ukzCcOb2lGi9G6L9Rt7lYP863m2u0JameOJs3
Ld/sIQSIxVLhQo4z7zokPrTkaenpCUst13i7QmYPhg1uWLbPQP0wv8Ol7vBW9U2eC//I6RyNx9ZV
RnpJ9hjolUUyz4dgz/s+pXhITeZj+mXFaOx6Vg+qkTWnbmtJsQcgV6XyLXVk66vsK2kUXN68wOmt
UsMK6vGWd/S4R3MvqRqISpzXiMnNP5UjCRGAMBlXsAYAdWei066ziKyggEHVEZnbUOPITQcqEW7o
lHfCdGHm0tzCNukiiiLbk/2GBifAhBOTNaaDR40U2hTDuOHzT8a0UZ8+cktDLKm1U+dQfqimmkrL
WGftia0sWhlNVjLFe9ZUIIzaTvkEESRTaZKfSFuufgHDFII6EkWc0qSD+WhX7s+dCi3fzFEZxXJD
RqibVpLX3YIlC5qv1z+Nxyggwtm8m9T1cdRFlEKbionM8OSrwKVgNFHNaNugx5dfIBEggdfwaUne
U2Z0Wcffme9QtxTGINluoTtkK5++daPRF8IfXWfJEZiHJ0DPj1w2uTJKWCQ3rQBgw4d1eZCgFPlJ
Uu/dxszGPy3kXv5kYCyXlciijFI5qFWiOCOEsRPsh0NvOHAQVGfc6SxqBgfA8NmZTAv3161xwNAv
ZBDuABlSBZabJI49bkgbp0DR3zVuKMrxWRVyDc/1aXV/IsOd2RRBEHNZbP78kzrVHdeBC9r/ljuu
ef9ZV6yLSk1diuLef2pYpgsGZ4ojC21JCj9Y2s8yOOtqaTTi7MWlxHGYA7T8v64b+XTsZTYgj12J
v7VBG4zSXZWWfRPdDfjLwYJZ6TAlMBhdkhsG0NdOrfUet/VNWmUdbKGU0//cmX60iLMHufi+12ma
pZfk6wFIS6FUW1YdOYVpgbhndn7MNWdJtuKG0ir6ENeBosS1tomLUQOmJdaEaxKekqyLxxlRC/6D
dFotuZDvEb6iPnYP8UqjiQuItsPsLNISPDRqX5kujA0BsgOl8kFmBCmWfkoMz1dCgsb038HsmR48
ZBEVW+m0PqOUzRJr5fvztqs7VkmlU7ICxt6qUQybmsQTUhxoaiyafpA4p68KhYpMyQjn94uobOoP
Lhj5GY8NO18c/n2kl+Sl2i3wRk+iE+scuxNTIFMJnGehkYc1Dv1fN3xKYcPVOl9IbCtkqBDKFfGY
i6BUH5uDtKkM89ZPgkFv9rBkauzsxagMtBO6CYrHyul4DkTP1R/SPzviKCxP9qNwvg0Zm+FbMFtZ
CQwAgpQNV4evjaPPl9lDnfiuK9J2jjVBv0MSvARysJ5RQLtj7UBEKMUYVO9SQvHmqLZ9mHPjXYa/
k1v4VedyesXP7CRdhpx/QEQPi/OpIhaYc4Jz/vII6dzlzI884tCHbBbYZ3B8ZYSIp7VqnPtx83UL
74D/33KCueUKbs/RNS+0MMOIJ3Rt7Ok+XAH84zwqaaz9QL3nejRE5VmnVoNis7uSO1Oy96xhUu0L
ZBBTSxBep9wFwXZdZH2b0Yx9EEc5ODqLqDwtenIUW+Hlbp0KnpEhkBdY90ziaw8CQotYKE//7tv0
lm6H9/fjdSKm5j28MZWMnix7qbooeRpz9ZrY56zkep0apLYYkVhgabC0tQ1r18Kcd2TYTiJ9T4bu
LE9wD1pouKd6NZGG5o8MJfgr4cKTNkG825UCxjohS0fB0DezNtBpIIHiPfzHMO51tT0kEwoGVkje
JaryhON4FOYOTTrmKWGb5F8h62BrOnma8aouNpSYNbG5srpx+xPLwclWF8AMFnsbjzrB8Y0MW4yy
uo4B5oSqfam/kYUwD7bKEaybyeIw1fQprSUej12U52/VRHEyTwMXQP8Nawq6mUIVKLMB/Q103xjA
rfrmGMZT4kK9VWx5natBUzHP6K21FPuai5QChiXgWB7ddCcXtUlauBO4ouSamkXHZG/R4kXn6slh
vUT6pEcYvb0Xqx30C1JlEOn+1Tmg9HtUCitCXuDb1JSuxf9W5rJS4JciCcHovH3okYO4FMPIy2BN
ZJeYqMr7tD0Q7VN7nGaWUugGXaK3zGn7QVgpl2VAuoBk1IMiWJp9lrfIe2pVDsB/2iLWHd+2WqTH
/jSxmwkSzntInDFi4LFdNnweTpDS0tRRVHskYix5GwwX3FUnnNKkpHJlhf214ZsBgIzkXcgzdbaL
fZxbJKIszNQ6wrSkbzZZ38FL95gK+Q5wjGgB6WVIS4aUuHRpVOTiVwN1kywQ4oC+iii+tvVGu19+
dxh/o4tWH3GPaB7M+z7Fe9wlueSsjBlM4X6e6EojKVQVCWp7d36Gae30MBArH3oe9REM1AN5oCjJ
l5H3OJWVMCxjYgMn28nDWANfPbzK97xzGHoTLeermTcJuIl3iGyB8dLknAnBoFrf/qzKGXaKzK5V
+Xstt7ibGviEjeWvunz5It4b3bV3Nwnl/vtsUhGU/+OxE2mfiUP1NhyUWWTXTN65BvF8vHg8fV8R
LWUcN8KYIrMWgvVgtNSxAEs4zpeSKC2VWmHPuB3ggzTFbTgBcttX91kZogJzCYiU7yx4+6QEtW25
oNaYS5jJvUgZQhGrEqRuHq3Z2roHwbToXQ/FwtQu0Q/ONDPyVzHX0VrZzEP4Wt611H7YrFUnQvRH
e3ha6NPSuJkocauW0O1DOP9XbkCGr4Q7pLL5/1IoTxGv/7Q1o5vzBLvkcu4LobyC/rT62WSk+JrK
W371V4t6JqQFaCspgrFFLvxGXfgdyuFTZ45v7+6o3VWm8YGFZ5OKrfTDZ3YwSRR7aPVczuk4G18p
tsWugjT3lGJ74IX0GiB0EdKv7dg2BNqVB7rQvjw2migM5+5ARPsWaseFj9txBhEuWbCj89/uA5F9
wbihImRsL2SD3mOHWPrM0U6CbLJWaZZLeEdMWc29ZXDz/sG+Amm62vJetyw8hZ0Rvbftuiqo5YWu
SZMtSivL2MWhyTZ1mzJU5K6XGRMolHVeCijvfAgJ+MlTucfCPUH4h2bGTUoT27g5GXSZeRhvEkPt
1gvbwq7YrTXPvUIs9aXhcmgCOTPsAbcLagRsdg4VEGkSABdAG2J75oZB08TKM8HywIiy3urnqNu+
taRpYPIaJDsdFP1clyrWybAdZ/S8ZmIhe+i4ikqcnzS03VTfPmA9HASdph7QpakSCIQ6SsMpOQn5
crsj+yhljqU/41hDgaCXM9HbatEJXLaygw7TgF3/tlqi3eixZ5ipI+q1gdhDcT+5oOG98DjsW1d8
qz6xzSpxihBkz8B/edi/NP4yYPhWP/Sv29sP7UWRmlzpt9Dhv0kQRqG1+mKV3RvMMgwyjiQkLTql
gDs2807idyVD7+gAbczmwHd9lmia9ZjSOwF29YXpFooXdZ2aZB5uaELKoYOY1/y89Kx+hvSrGKkg
kmBTIl2wS8vUEmx6v56TOPBVE3vBf5OzS2inrWu1Oo/G/7GpHWIgLXAhl7CxHCHzMh2an6fa8Kz9
x8LmA4a6Sx8/AWp/rwLL3PKoizWKBdANg8vYNrhi2pfcMdsQiwpwQ69CJTd1we2zlVHw/kP8IGoh
7BNLKi6jYqjtNsNTT3dPIuR1YxSA5UxaJShOrE0aiJ8ZOcifdb9aWgUraPCHS1BjXwgxhnZ0RVOH
ogttJNGUnnkWyNaDgKWWdjEBrOfYapW09Ru2e0vnVYrsA9K3enF/rUuQFIi8Jy7VTvA5mcTkP9Cv
SPxNuGyeiLA49+u3U5ntQPCzE3d2ZwmCcgbDGUTOmGpTapIp3FAAIbOf81ULQ+u2K36a1MllST/F
ErXGLttqDvtNBe+wjL0oG1TZhQzaIDQPsjbApYMQUHwdEmovikcxvRBUpRHXS/LDxgXawFz+hN4A
NJf5QOWRIiTuzlC7H9ENuXNElAzTicJnsZwMmSW5nVPZbZgrUk3egPjIckEYFthq/I+UOYsvnlVA
1+78TCKL1KpMc15EBS8ldnGYyE0aC71rAXpE2XTzEOPjhwwXk1KCPeBZi6Bw2ng3cmMB/0zuiRzc
MethI40k2u58GCnNrU9Zwl/KFpAOMfIzMGRuLlxknyE40kzEkyi3Opd1nJH/7XI8OT/321FEtYh1
lxnK+bM6YmmckkWn2fm5D5+uaLdfFQD2L9TsKB4X8dkr2jV/DOcIormMcooPNOgPKad0ODNjqKZY
x7Yd14vLP1sFd3yNR0OVtF8sadT8Txh1pibRFX7o2hnrch0ZrvLH8nY0F2iDtcrrGZf78eDNB6HV
sq6HHUObAZ3tD3CYRdsAXoaJlEQkVwG/sH7MQDewMpFDEwgIJLgTgDiJRzmA8/GLQZOt8koI/EgN
PIjmJ6wHHLK0J8Ip+wx5xq3CxK7avlm7gldNTTmNydr/3oF/6MaW06APmgP/ZjLuUyEtuOMOOd90
qL8kp4IGzGc6Njn1Xt8Gr9iH3K6iOvfaprnyfIcvJU2pEji/e3nLyh0aOX7wecNrT/pCmYKpy9b0
Asyy6SWkw8Zezal0LzwQibJnlV5c/FmYMOaGftS7xRnUtkDN9a8H/er4KLchBMkkiEzlunviks6h
Y/MF4/l/45cmtNkjPZcMGXTRV0NqwT6gxMAt1X0iNAhck6C3y0LMRxWMkVi85rGd7ndHJTJ01m39
Oap+BVXu2dTDSPDD43nU9gS1cNzzo2GWRL1nyR1hmBtDslPxNEoe01lwzQlILjiEkSnZoH1RAZz9
ZEkCwV56DaQmIyCZek3g8WPQu06HEVWvCxhwZYWGQtvaeZxOHopTITesmXKCYyWArtfWTsRVUkg6
nIWSBeBJiigMsLHielDD6+ouM42M4rb9F1ZxolAI0R6NZW3IE8iTfWrXihsFUf5gVamaQ67W23Zu
6gamOZsJGZrlVo1x/5wefgGVUmanD3daonzV0UyKsig9y9HC3NDOFpQA7v34eb9756mSv7v9QOvO
HECgg0WNznQaVXAUJORxnp1J/YFRhACSzGl89M1uCMy9TUlHIFfwB78ErEMr0ACZjCT7l5kHZWIA
Xt/mXgACmjdVotZ5HckG8vnXQzN16LMvqwAuRKto2/Axs8tyoF8ZbfU0oJCuBvZcSzMSj6R50SXd
tUpUlOQB+lFtzmzK0gLb+9ywEZYdiiKu5Ga7luo5qzrf0o1A3UEU35PTQY1w71iWNVMP9bsKOASt
YFttUbKOk1iUOGnpHPgiFCLLibrVKv5hGIqqxKzXLiEjOVkvnHs5vtaM25I9nrja1Uv8uEs/56Ch
H1m+MXXjNFKqCtqSi2Y16dvHltCR7JkG1t8JgQMnbkDGq4OojlwS37+RnI5qLMaQDK+3Cu1Bf7Va
eZKwWi18QpfnoQLp/zXDlDnxRi/ZMDaaXrpiQT+if9NP2jSIhPg5IzMczcK/LxVuaGmEk8gAtKX7
VVjJfgFODT/iM9SDW0V3OidpopF6XxajNoy9F90HpYGVr56ViP9h0Q8WF+QNCzS1F1CUoUfKswFE
UXKf85DzhHtyMHOv0UnH2XJx2GdQPJwbzhrXU7AjnZGg1C0nJWD/8SUy20Bz+y5Nqn7W3qBMuDvD
SmopGi9VeBD/HpZ8q9J6vQjV6Pt0/PLeNjBj+XyxRqfn61+/Pyw9Rje0WUJW5rOp2GHshU4AuZJ1
szL1ctKjWo2bDoBmqEymOjpclrnhe4+/ty+QHakLL9hLrW518xihJS+db2/NretGaCs25D+4R4LO
PGfHI6Z2EpjxdjA6x4TmfMHLp+tRlV8PpzXUnJrBvR7w81Kmvtce1z8C4iIINwTMPem91n6U9fhl
ahK0ypN+wnbzoCZh+kTVVjJwt7jwxZh7DF1SUbAjUlf1NSeFxIgpXXDojYtSOCmgz+bX0DjAuDBw
PPk9bNa2lh3yA3g11lneTp1x0AOKUmyHoKeSdAU9/fLAZIzTtNNCfqO+kCBHKpoACFzH+qxDl+tY
QQaFuqQpt4PmL0ydlhFg1Hm0cGs71PvKFRs8RJMvSu8dNMe4ShtZiMLhmVWmAtR62XkSHuMRLDL6
ES1tnaZdICJRCWujdovTsVp3I61xrZBln2+XStCrR1MP3PZ/QocLPsUdqTBcykC5cB2BqkQ2TowU
5bDo1tVSIb+bdvpkITgU47qQppQpaaOulQTP2bBGg36OMkehr1O9XbBOOJmd6vxBqrvLb0V9TXnQ
ksauyFlGPokvL9LFg/DA2g1O/MzpdEr2/AfIskm6uc3ItY8lbSTDe/5DMc8F/2bZLzXTgIutljzf
ZKDC/p1osR5R8ENQTTD3mrqZ6rHEvkJ+TyR5UmXOaH1MmkOeX0E89sfT/7GvXzBcOVgq+h3PYh7T
RbPtRzQEv5LHecEI87Djy0JI4LQ6WazvO/ZfT46+//wlM2H15j6UD4DFkcUK7sD4Ewvy01vZdmKz
fYMloKIsay+9fXCwswslq1oUMXfoFbPrJbiZDow+H7Tyd+LGyszHtcHqdj7ZOKPPgjik8bnCFmtd
vkT5MjyoxP3nz+oI+tULGHIBq/yf+V/j8mmnZKo86atfVC8qLLPiCohVNjuU3eg0TW/2xaRfxd8v
KACF5QxpB0z2+tsFGRYD9z/xapppgXM2t2KhumdxjvsI1MN6TWpTsHqoEAac+NyQ8d5ia5a+w+mJ
0+/eFAPYjIDMPU4JTVbX/P9RAd4POiFq2HPuwg3EGZwJuJg2SKkCNlN+vcjIOv4HnJDFMlNWW8H2
w2FQFBCUK0MSBJ9mEQHNupNN377By9/qDHLwUgWhQ2BViicyZwC/2UifruUz/B7nijvOv8RNNyXo
laRUe3hHqtryswIraK9wX+KNF1onUSenvG+zXMpFl3dIsSIDFPn8qBNcIoSnDZSi7KiL/er2CqY3
NzykzoI3NKteUxvLYFhGkqTd8VpNRf/glj++SRc6CJd0PaBZzM5RBoBDdwrXEVAgFelcD9FioUvD
S5tO2YtcXX0pA0fezJA5V8NP98DYh1mDrLUIpXMpGC9m9f8Lleg3OeCzDDOrzqaUcLhiI+PWdtdR
S6U+04MCkVX4NGXwI9lfpWlb2x1YDQmpIpKxPfdt2m9SvpJgSrsoZDnsW5zGteSVZLZB6U6IdzVm
btz9MT6RxednGNcz52KWK9HNPGJJ1KXbh53bYHzIo48vojvjB+IfBQyXhnjb62ahVaHU/4A8cOtw
QkHAn4DBWcqAU1RYnwrCd48vBlbsj7CWffxvE36mmXdqC1dP5sm9Qv9amxV0nR4UcVmH44fw8976
YAqVZh1MkD5oXRBu23z4QikQh6J2CnGOXnWFnFtleoq/bz6o169uJwFAethKLjWJZivckiP2+fM/
HhJFWq+XW2ZhrHp76ZxbyzaMOo8d5XZtryj+v9xfjvALzbcw51GHVrBQsJW69L3i6BoNO8EGFTpW
4nN25J8ONeiBkdscJerWuiAElHvDSWWVyu0IO/Jgc07luldjWza5NXXXiCjyLZy/2L8SYrceRPdV
fy5NwtoxysoBEqgjYr+DJ5I95uedkO+rHjUB5HousMLBH8LW81sviNVWqBHQljjfyoeVSquvB+jE
ASr0TZZ7rr9qFJpqWMrFEpZgjFq+LJdma1g1IGjAU8bEY6KUvSomMDBiikl4fNUa039GVTsAsO/q
rURr3r0bVJx9KU6TrtkLrDXJKKpIcdAnhJ5Sh6AgkWGfUFw1kZRBloMNOgFKCDrwiR+DYUV8QyK7
Ymlf8TidahqPHHMYK4EayVH5ur+BqX+35gjglnwn25D2F8f17jNkfUCQ3jeoOFPu4vVOen3dyYwz
Nplr0pe1nPBtMziI7ujZ3COjrlXcXaEDvrfZSdkLDNXFxipGbsDpQ/XYc0nTgvptQ21VZMYoIvcI
SvMxhHKiUWbTrRvUbgdPRcP0YC+g08+Zg7qSdy+ZEfoTTP9wLGGQtftNd77stPvsnHudSE/oXvYr
YTOlKztBfSAUKwEmkydcUgcbnv2LxsuAV/z58y57xpHMnogcAfYSEiHE9ROle4iQ6dLqMFx3X8xc
aNig1QTgugre60YBGwFv1wQGT+NKGafO8HLrkyHdfmVJvUj2r2+hy7HLJ1uy6axcjaCcvypcgfth
Jc5YG1007YE0IbtFwAdlg1OX4zYCH5umpE55MCjKfbPPmbCgbeMBdy8CF1g5sDqB9b6/1mrGtx9+
MGJ3Rl/2yCCrVZdZo4L/JFisCkt0XamynDVP5fko5/2c8HpL6vGnQ3+0oNs4KuBs5m2J7c8vCvJ8
B7VZjxbKm75dtTLzUafShjkVfEEZNELt6/eRCpQre/N5MWfmTYrAc+flZCCs34bzXSAc5XFzX7bC
HkRXRyfwRYHeo4oEaO+9R1GE7nGIG8u/vosuPhvR+geNJqu39vCiZQOcR4yGdduSM5uJDXn91lXv
Gzgu8RzUcxcnzwNaJcqxXEv5h4REWsYMVxYM+5a/FRFLwGSBR460rhZ83dqltTUtC1B4B2aEb7sQ
dlfVAGKNSUKy5CjI/0+of1WCpCK9YMTBASGLCmuPElhsv/C5uEiEuV7TYWwO/BOrvOS+cqvpblBK
BP4gtLBC5nb+MKO45dW4yhCgKeFcktYY413IVFpppbaepGlp9QX95xn+tU7eSrPMCE3F0e5Ue0aF
OK2swXTYVs1767vnuJMeSHUpO7rUdmPSkAXm+SIWJ3+F+g1/HyCmZhTIxNmf9+soU2J3dnlT34Je
yUYXWZR9NDpyyT+r6y7Gz+A3CJNs0+bhri/xjUFJ+oFtWLdI/xtA+iUf2TXzFWVK/D2HUI7HDPU7
x5P4DAX8egoPquP1XV//rhp8VZ14/8PCK17c5QvX8s5URJwDft0aCI9vlE3xJMPzZ6ige7bayF6r
3+T0ln5nn1WSNBWCPORuluYUx1Qad2jsuWlThqoPWQXOav8+TquMxngEXDHhKcaUFuxuvMdMWm94
72R+qPHfY6ruqa30hvzK6d24tIPHHhVfl9sXA/wFx93Gm1Stj6AI6/CxqCtR6+n+DIcWwQ9622Yi
J0JzgxCK6tDbjaxzAv1Am3E5o3Q5zu8zWzrxTQUdIhoZPduWTrMZWQO57hgjxXodp7JT9vRxb5xm
jpj+al9TDZzYCU8BTO4vK6/oW7krR8uEnR+wZI1XVP+SxhenAJYnY/YCfTEG2xsAo/OgNcUnOcOS
LLsOpf7s1yWFuZnul4Jy1D+DIwruwC5AbJcAUDP+1wDs823BSvctSxFAvRsu9Qqjxcho0boa1Sd4
ZPafagm2uEjiBvL6D6SVKu6vAKNN2gDZpFDXaznwwKWiwiy4xHKHhDQBS7EqFJGw1hDT8aMgAtRl
JsuLm1Z0LJCuzpR5djN/Zjs9cIXN0vtZhWIKbhuQSoW2krLsPUTXIDfOMRW68kDpCY0Hpg59ATdh
TYn28PkjwYLXWHpVld8IaBgj9ugwTJWghGSNkyqbc3crtdzg5LS0yPYW0WSbR3qRAw9KYMX1eXmc
e7yfD7xSU7JsGj49lXsyOj0uY5sOrlWIwxyYTfP7dZX9F30rXdHmvatGdp6pd/1ocRCt5fuAemWT
yCaA125C0nVNSiUqPsCIPd/kh0/MkgPT5yZAeZcugpJan7bDUBGN9szSS9B1c6m2UZjsrnX15O5E
ujpyuMqVqbOOjXH1mExs1nvZ/T1nXm+C3luf26hlE8bzb/pr5D6LNL2gnCZsZSHW8oM+Wcv1k8lg
EOZKyR5pIMf9xw+cRPHlxgKbvbnkQ/B4Lyu2FezLmmZyqirZPD4APtjyvC/rIn+r2dl2ZiFW1C6P
QxlebzztG8d/RN4nxOMKQggGKRp90dz7lwvKQVng2G+acJh95vqdufVB26wpwloEqlBJg3UBMWvw
UKj8mfp7D5FOXzg7utvUFokYtcLezryhfZcS0ZQxOetaNDTqWknOxC73vDetOII69BYPtO5zAPz3
Zlvv7z9GsoiLrAABu82cYDT/rO70elKQJNEs+UiwRjTH0CyvKxYuyTwK678/ReZ6tJdxcJ0G6xkb
FkkvhyjekbYxzpikFVjZiru3utLmgbbdHmcE6qFTzXrKkYmqxKLYk/sZErr221xyndNhCbVfCtax
Sw1Xaj3yiWjWGYbxYSxJ9NFwiC/fxDcqtLrslx6YO2AV2G/K7vKwXfqUO7WOg6OffYpSK+X5BlzR
ubwOVosZLgiNX0SNiYB6/OuFYiWUlEDgBkKnmMm35+RaOywWfKt7Vethc8/KilMUe9A1pdosc9TP
/h44P5XIdzi6ysVFiV0a2ccqNw8MMHs84h2hsuutz3p+cousgaygV/hQuKU0GYNfei5FtfF6tipQ
YiqUgCV6w84yowteGv0/CkZlO8EBru26YkrqA6wbGkQRfChqIDck2IZwtgx91K8dS+Y68Zy35P8D
k/z3KM5KVZF3a2cB/0QWjVbilSTflSaab/N6hMLfqPW4odAxAg5KZPq718361KcOGg+4ZVoSfmY3
DmQkiF+ZMdasFVzE+30E+Rcoy0FgQy7ski5Y2tkCVKv4+j24GXOk/0UeKeVLKC5mRhzFkIZucEq4
Eqn/V0c2k/31WR2k+SaPXHSZVe3q5M0Lj7OXdhBwa0uVOq7Y0e8jDYyrAZdCrkhSlrjDmPSFxm4k
HLOdtdgXKHEga9Gz19AxjpjdtdGt6PDMsIhxmQdteqwMi0pjb+nQeTwTjVXBfD68GGYUUxH0X2+4
ilDcK/yeyol/cKYsUNFOJ5RTHUCbPQ0mQxEU+Bn81QOEnnpcmiiHf8TWaBCh1UbUF6Bcgg7bBN+j
6myTTVFVw96N2PdIT5bWoKZlY96CW+6gOmLg9+aS730zDLLfgCIXLOIHcslpgE2vfKBPYp9Dj+LD
pvb2ieMQMPlm2Q9OBu8QJLgu9byuESiY5zRL3X5eTUQan2xR7C3u3JcArnC/VedIRcYU390Z3NCM
NZ1tUuKZxjxFt6+G7dtThP+s18igLhPK+4tPuqO5GZSsK+xpBCAD5r3TIsRWjEJdD1hpD29D1nqg
+3OHbqKH8TASmTHRzdGO6UV5e5cnDtsyvfHgd3/A7a+99+LpFQbLq0G11J3ud+JGUVcHD8N9e85A
ObIzskdOr3MvQOqNSjxdw+812y6vBlOtTMB80PH1O1sHE+OQtc/AOWdI8gVvjIvhVmJiNuaY4jeA
5sIxWBPB2FUmus9/eqHbLxMkg8fQVb18IjrJp6aHHEEBPFot5aZSmk0eI9GdyRYlptZD1ENCOqMY
YmLiUPhvWqIDJ7YxZlXQzLvwJuzO6msSc4O6Pz6mkNRzE8AwqC4mSdhsm7skzeBxN6VYmNAmKIwl
78HvI/KnDuwu5iDCpdD+0nD8FZ4dM8RopaxwKXKsAOhqAc/VfofZd661A1IwtQ3jVh3SM4xH7wLz
/aEbB2z3lK1Z7B8IErYCWz7q8l4H797QX0yTo9KfNMLNpbVLGn/j+SJysI1BYPw5WHkVJgcgWO9a
wkClxoAxRTUPl3SFT7x5FQjEMegKVWaMrt+ih21QjFHcvBSNvBAma9evyyZXPY6D8FtHVEWOJqVC
/oCjfQe4Rt8I6Jn2AHpbxQL1h1CncpFLq1ymqs1VYGxoOR0sTFVU8sOn5A+g79ZryjPT5KfFlMhm
6FStONWLWyOdy9fMHUXk3M9aynCnOYEEpT8yyVeRQHjY+yIdkkYiG4EmlrOJJer/mgBtGb8zTOjF
O9j1XikRcEX4tC+m5Qyhmg3bQYPiQqBplhpd79qDpwihUe0/vo9OvKTikt4XNWoKykHPMt+i+zUX
jrJkCqs4xU5wcyMjFTbPDrPwzqmHY7wJX8bCJzrWYQEhYOQgoe09oM9Rq6dJhgHJClTKxKI7Gc11
Jl79DID+4lSPlMmCIr56CVJV5GZ7u9HiM9Pk5LiThzUhJW16ibZbwXa5cwqUm3QwFIWMSECwXshQ
Bij3l9k+t0pDQ9CUZjGj29XHFJ/qageq38ZDsxYsinnsiiBSl+OZ1FVd7pD5jXJVfDS2ln+tx6Fn
X4BRnh17WdwDv7f6I7uZJ02w6mU3wC7WJNiInpLpc8wkhVcq03RDj0Mly6ZuudbGjHwus3kL4u3I
dUhfYCLV5w4idzUUs77TwJ5s/Hz6LV096M3BnJfFS3VaqHtFUvtTvZ6KJ+wC3cAX37dqAg33NYj0
3oCGHy3Zs/smpC/NYsiXXJv+CX9UQFk7/aM9ro14h9aF6+hwE6nV//PGFUCTpUNdik+X0rVwg3EE
a/Ap+PrjciQ5Wv5IvatpUHfEJvBdfNcM0S46cNcKL718vYeK8BFRSnv1Beu7MOo7nzZIMUfFdjRv
UZSZQPFDnMZ/LTduA6HScGyPL+nFfdz1o7aS5oqdcl/H7dWxkUnbMZ/K21h6vB4AxS30l9n4B+iY
/pTcmrCn77nD+u/K13c6rkevxXX8sFRTJndxzrebiChSESUm3ErpLC1JDqfoMUqhaZb0Sz5zf9SQ
VLFS3RT+CVgd1eXv9TFaKzOPhjZ8Y96qX3Ql2eSf4GcOqJtGRJgmrkRXxHYT08j/nLFJc/veCivl
4N558kag3yqxVm1u2gKaYMEhCeNHrIwOMTedS/Ko0hn7UHYzWThziWZewyUhVvarQP05e9FBdSet
IPb8SotSpnsMIkpDHgKack1GBJTAFh5d7oEpUVq0KzMjB2t3Xz3azUHb5YMDAwkSdc0FZUNRYSJJ
eQxfY3HKfZ3SJ7fVHqwsMlLvRBMQEQUeYNxp5XPu8Y8iYr5eE1C30ghVTQtWjTFeq2i84CCwrvZD
hnNW/bewigSSmO+6krriUN0jUV7DG6r0lReoHLlFUY3Oqx317/+aPsHT+2XZD6s4QeI/dMFuJlIG
z1akz3FsqbYv4VhPqmIlxOIU65e7Mvo8TxQp/D08bxR1NmCEsEp0Q2SI1TOhvDjfG9Zlgp/mPQKf
ClPqZF7MLRoq+FI7NBwODcV6kl8PQJz47dBRmxaC2aN2v/i0eMtip/sE0sGMMahAA6WWBSfdbJco
lkW+X5YFE+05DfY5Y4VcaVdhb6bcZQKTRBy7fVhnx9gsntj8iyHu9HJQVqeeusdhHk7L0fQA4taA
wEkBfB4+1QrXH9H4aYo/qzrkJo7DFYfc6z3CqOV5Mq5TuoSoB8KdaSRLThBPqSpTYzyYus+5MIdV
00uWSwpZMIPCbDvTriu9FybtH+cARIrPoph7ErLZKpGnDxs03EHhVa4K8R0i+wdNe3bHq4YGZoON
XVTqXyC9XIWAVPOT7wnpQFVf/dME6OcnN5JwPTs4Lk1zeEinH8DMtr7aQ22etHaPkloklPGLo++6
1igEenEeWM6D59rM+YPRIsuDo9XYyQ7GifLOAi7UFxkUY0hRZ0JU/VEo4fJHdkQS802Ba3u5P5dM
hrS43DCX08NPiS8S/BG0Ts4LW0imeUY8DinxIOQ9mwLEmVMskq7s5Sr/qCTb+jsIBe0yp5ifgJTZ
/5HlZMkEG28DBG6rFu9ko+lt9riVTkZsfPVRTkEjqdqR3dv+qKkKhhIJK8qgcrZx4hbBgWRK3VoU
35WM1o6X5FWtVJNcP7cjgIcgahq2wdcn6Ir94duvSgTdwM3IltVojNR2tZNE0/qmz04ZaufIhBR3
acWIDozQ2WCHRyCZaD1rOdjU2E51m9QNg15DbRzlDLkjEi8ZmAB5rWHtbTVJ6+djAKwbxQZmBRFd
vEY+xkwNfXS8GeP7Ywg97OfkWpXFh6+MNJ2c3P9UCPYNP9WekXD66PkNwnIQy0s6SmogRoL7SeOt
ZkuCJWcCdV121T2ERzw6B5tOvg0Dnmb/bW67w49Jq78NRNTVhHI/6PEvwe2FEp2kSDj5fURFOBBU
dsTLHB06FmICiE+2vwlkEe1WRfI1KQFoydgjqRpaE52OI1OFgHhRDwM0XbrA0LMycAaEZ5fwAmyu
UtREYX08WqMQ7Qad9OdGWe6d1JgrrTdD/o6yAZmAbcF/QXW7/12LexTMZDESq9KGLyfo5+k3fOkK
wuTGb53yBkjbQ+etU/koKLUczgdBsppU8jjotm6R0BBTYrdNxeo2qlQdm+7DKlVRJlnPQTli5Bvd
oMWu3QVyL4bqTocPhIFkMb7rAMe98dPb+4utCvLkzzULgP6OWJRsWJeS7gUJkwrRlBZfKgvleOMu
JvKgAt1C52tf11yd/cVe35SrsHnsXAdMGcn9rwnkDBdSGl9FIQsXIc4UjQBiq+KoS1oJ4ALcJIkN
pgoZkKLXtedjwt0R4EPFkjNG5GzvqPeV9CwDd0E+WmgU46RBITvOk8/Lc0oJ0G+A2PV9InicXfPp
4xvuCbfv7lfmtx4PwJEUMOgcbYPfBgqsH8zfmzbnBUHt+0NF8t/+wg/oVQit1UHQaj4sRLL8hBR1
T1Juw32SLH8y355STlkUNqixZSmpgVwjLZoo7a0iHn8nh88KeDwvmSSFR+sYXPNA49+Mp4yPb95S
UzKLEj5TqMazS7h+xzft+CPD4waD7GPrRcg9nEdqBaNBfXUU0JYbUHl6iIjk2Ld0KBTmRlR7FYID
v4IF+VNPAc45lzYMyWopOYsOdHjh+Y4dmEY9h1/j35N7cal4O7YBKapfh3jq7kuKe/R3TAxfzytw
C55hG14AnoNwLwQgtkt7hoeXgdDSd2nzjN3+UrZdA/SODlG6B/ezmu+PMzq2OLldIVlVv36hBM19
BnBQpD67BbuEKEji9wDFa5IRU+81MCuH8wHCGDzB8yWanb/noREs9KOHA79yeIErxVShUcqTyCDO
42x8iKAYseQFsMJZoq09V3tRR2PKxFGwbaLdgklamQwGwls4cHJ72Wd7QhgHFvq7OLDs42aw87hK
5Ss/W8oCdnp2dJVgmwAtl9WWFsVDdgLJ8q3OO898B3CVCAmxKeF0V431VyNWuXAHUFxsQpwHgnS+
qMZ969wGcYLDxYUXl7GkSe+DtfHrDk1Ym7m4jSPBaCkArBMoj0LtBIgKDCuhAM2giIh06cBRvKxb
HO2q4u8+xCrVkMU/qrEpWp44/QBtXkf1viegvzP6FMe2VRgpyfgG3oZsgy2e5dHCy+GqHq2cWlFU
1uz8V/9biC/2qgwbCLJxc6PnXrUcJFgnZiMza1nbQqi0uY/5vHkM/epFb8Ecufq1oXAT/3TgymxZ
+diqkL6IrgHZBpyNKHkBdG6zPoaEQjgumxQKiP9HnPj3IA6OmyXvh5afr62RXeFZh0KpAWzQIZbt
0Ue52ZvVNsMgbMQaxPBWsKv3hbuQOUoBsO77W/wh9fa2SL/F7CmYpNUWzEvAG7edpsnWOU59hrsa
3sbX76QC83Xgd8ZGEOz422FORWI2HEpC99bVAggxhiU+FUtxKKpVDsipKJpolvSJBg+FBD78RXYd
o2vSVPg8fgqPjaJ4WR0NPD2sLCygHNDCKgqlI/hLcy0HMHNV2RSxjVO7yKo6yRQ/3lmS0UheCWL7
UTengcg7kM/4vPRJc9auw6ocjiLzL04tmYbpyDIciBgJduyDDc20rToy9dZF3oWPDUJa4IO9eOzv
v7NGURugrNXSOgcPNmGedTVHCA670iZwLNpSGQp5dqZfcn0VEY/2Dk29PwyoCBxN00m9EUMhnBhh
xD87jHaMIpj9aScj44SG+c1iBlJVa9Dn2FOBk6VLGD4SZI0rroJGv3orlaWV6teuTc62c4rvVSsi
Hy28IBzDvFzOPW7mhYGKeiWH/rEbr7jxTMozZwECC021lzruZZKoh4BXeqGEzvpMl6Us10UmRKIe
1crjlUFWGTawmWXmtTaLnVo0ZioOdtQAN38Z8w6SOoJbaDgq00d2s3ClJkRgRkljNZzFpc5GJKQP
BSs+mSryyiGwa8qN/TIpB5CfXUT2IQcdPZrAoNAtEFWD4GgGkZp+OO6r0XHOFDhfxdlLzSyuJ4D+
9oiQqZW1AHjfyYEbQqMAZD6rwAWjVkcRt4/3P1EMStI7G9lmso2pj2yVOoV0g13KQH+eN1Scri1t
cBdevCx5FYncMuhwlg3ZWVcb3Hs+akSKH3FkuKsQP8u40JtVcd5v9fozffguo/X0VFE+Rj1uce02
Hrczti8QfaT7J4wtRx7WZXqxKn0Yh9D88xGGJKp6A8LiwofVb8j7hMTqvHa4ih+ssGyIvdv5DrEg
bKWgS1QrJHA1BdXzvi2xuq5C4GlCeCJhmOMJ+HArpAm3hL0msn6k9XJ2hs2YQTycd5Zq53rqss+p
Gkl9urZW+59uqiSgIfje6drM6yULiY8wGvrQzKg6fH/JXT0iH8Bs8YbLsXSjjbXIIRhGsPfxZjsz
t6zw34d82tjBy+p3kLRwO7qtHxMeedyd4qlFm7DNDB258LWBqKXzRw+x1un9XOuoLGWlKKsfT954
+JP+gDt0+oGS7KC/fE65aL4dhP84BkY6K403sJ9SpEwSo2/G4IeBdC/OF6byn9Y/Z998XrBVN8ww
4CNunfqOpDPNevzd+wtirXGnRD1PXqaXGbfykc6m5NgABQOQsc+Sx4B/lB+ttM5GfKD7eZ15hDCt
Vp9VqXgnrXpynkp1CBJn8UPl0az7sSESvA8IJmFEI144xnfg9ijs9biyzG+MikXMfTuczBasIdG+
IEPp2dCApcPHHpZKj6l+kXPiHikNGGwyx+BizRW3wbJ4US8csBVZo1NIaeL6liC8d1jYfDX+WGNX
zPtWJgA1SQjBisf2aeXUtYvLe+E7UELiU4fvI8MMepWoPYV14JZe6MX642Bdqi6ERl2XGB07/76S
GW2zMab2T0ZEe6sv+33YBdvc+39ywNBUNtDzQVbyORE6Zjl7/H8EkiFhTH7GeShlCBpjtGjLXLXO
2/wkV7JUYGffaFKY44//drFnF8KOHdMPkinadE5VLcr2Eaw63vBwi8il6NXVFVuJ4LOVV0l/jJWc
qSiIcSFEqRAt6xHAyXNeCHRpx4pc9legp81mKWJboaeVifSM7NLJ1bLUaqXv2aBgnirPg1prHyDT
vbY8TerfSnRyNyEzrqQU0Hb4x/UREiwB6L2LD7b2Cu8ISMkZXvFYSuN8ZgrroHeqCT4SGNm8mo46
bCEL+5A2bKrB3SWYpg5ZYj0WBEe8fL7zrnTQ24yAUzWVkcf36QyPIUfn2uETCb8Qs8HuXD1emNBJ
3XkpuRSFAlrpttdV1FexMB1tvq9iiM4Ui7K9A1ct/JaEyccWicD2Id0Ce0oaBT0A+oBh7xCH+ZdB
fTZCLsyDuBX7FtP/IPGtOUnrvd0697N8W7NeBWeVS9wKmttl14QjBiTFPR3vf3F8Tg+xeC4WBbuf
o9k+u1NLqQYz0jeLPZU87RWv1pPr9G8GWQnT92ARq1vD47/3RrQBhjzFrk8B5wmlumPzTGguYD1D
ISBzUFEEaUvYCs5GV5WjnRbZjlahWlWPv2HZktF/SUvAjDfjLO0bWn+ULe0+iY4rGKeRq4OLbo4f
Pqgyvuph3NyHRRh3884Td6D+3O0VhxfXn/Vf70wzEse3ftm8dlfUtuAyZ7pJiMU4+oIVrSHYWl46
lfgyqeBi+cNSz7rbn4foA442unNN0R+Vr6tYVGdg6Ho/ajyufdgRTO93/siWse5frpKsVo7WqKMc
Z9MDC+WJNeQ7k4kMEavab+t+v9J0pDEcOZbx82R8oneMjDdaQ4psUhSsmumuXJvNfaRmJXUQ+gWS
d4uWilMURLEyhNB2uMPo9BF3vjsv6rmCcTs83LOZ1cpiYtLkO1bQExirA8+gUKGIiUOy44iuoxLg
+4oE0UoDlpgRIREZFk8KCLGJPaZoLuPoN9hoeF2PYspky/dZtsD3uyMldqA4qvJpcCM2GjVf4gjS
w8pdy39A4/a14vGTf9a60ilAL3xRz0vm5RquVjiJA7cuBSYFgswadPC6HqT8W6jTJSN2nCz+Wy+a
Qv3wIg4cx7XesOO7IWwwuvKWlIKrjUpC5oaLitdiaaAPr8/syhHicldH/tOiMtQeDW6NB/EbLvJp
hUTkJ7f19lY4XAB/LjB3axq4g+Pfp7i6ZiPTOlB2F85bVRM7hOC5+SoLfBtULZS8+BowKkQlATP3
gTWDQKKW2q8XxYqQGw1c89preOnl8/aU2AHO/7f/2h3UZCOutrmvwK1CdhiblenBBtuKdqErp8l+
yCc+/UhkV3SnwO69EBgpem4JVO50OyW4fEL9Mshkx2I6aBn5aaBroTgPzmYUIXThcyCoTWFgpQK0
QsGo5oQnTeOVZVtsQIFLfAbIMmq+oI9Ao3u8t2MofimNSz95TuuQva9yn/jb1qJlu8CbDaq2Q3BC
NH0t9re0y3OhDCcjhsVyKHB5eJoTgV1pRkahhLMf3PAxZEe4G0w7jC5zsEhWuyfOOMRljD7dH59m
WnEq79Iklz9Vk8m20ibHkxZ0BJsxqKZW5TfrA6kGApSvARPP8G7x5Rh/wNT6756TWEPmYcrOCw6T
nx+ti9lQhE6X3SVn69eawQxXiWXJ+AuQef2zv+R3oQVq+ex3ApARRBbOO9Oz2//kx5qIb5GfsEM4
AvpR4WpppRKsklkyCMnaefGeB8HpcFvzQliTx/Pj7L9srfttsPYXuAV9DnZNBSHHr4lfiTDIbuys
REDjLnPycF9fAs6zGXUk2XFs493xUHZyOrKyHQXnYp0RTkKmdNFjKQAOTNrr1fvSpewFtodHAWDV
POb7Y/vCanFUZqpPBKpWNVefxhpusehU+M4b1YpBOM4TNjIl45bIbiAR/xFQlsTYAgVVh/VEm2dv
llGLV5U/9Y6swIUVY9bBuXJI2tkSGqMbj4w7zn8GjpXRkuCmj5xDTThJma4gVz3rRek+dW8rpfpH
uo0eQ6gfHXxy8MJoPy9B2S0hVbfUmGquCe7p/+REyw+3rl2UsKr3BuzuHeRls6AS++F2sDOc1S+i
KLdQ7fIsUQtUIAu7pvj8F8/HZtY8sVJKaf+7z20Y7nu5Z1jwR9My5wwLyxOhqhpvkKwrxXhnUH2s
8J9z7lTfta7oXMpVQ9ioLemb65fqnFzmwoXhEuCTYmQVkt3z/FL86Y5u1reRRUFKSEDdlv/co0JD
KG77Fy1Twku8KV9tjP+aAV2XlAW8zpFgUHNK4XBuUHZI8XMZG0XxXnzofV8Jl1KFR1Kz2GbwC1Yw
CKnbkoKr0yBy+jyd+XGYiW8jBm8bHpHY6EjB6Gw6U3BfEifu6hjiB2fowJ/4yP3pnaXo8iZaIfFb
HksF2fOQx2FCI4m0zAmRjqzjpk7DTneIY9xZDHGfIh24OdgxwlIwda9IyAUxup1ipINtRWZjh+kN
QLB7eOms6jIzy0hLE3P9A9N5zuxzXyOXMOUDA9zL1RqiKdk510W4vgeUbHTja2jYzA5UVa06U/ax
3LpEFYEbiQfaUY3zyAU0vMSWKdf06C48BGkNEgEyJvWR8k4td9zKn5Vr4Or5XXtU2KQboaL2oEiO
hQMKh+pN4fWwoUo+D17rrtyOJBj/7l4h/E/F2eLAeWNpmVQk9BvkWueSWG/1oCxICsRCLF2ZM0tO
8N1zfLGha8ckNRFJ4Aduq4xLSnlFwYm/xf6HDd7pLGpObE02DImPDX3WarsLqYem9D1BRRi7vRqu
NBYPF34G+zjil4P6CkRltgL4P3MkRinuHq/5SZwaLbFk0LR2rLHRwQJmnRLODqQmR5Lf8cbjE7w1
T+C81VnpJcIrDIiJ18VDx2K51KZcLdJ0pD0nCYv/BSTSVSgSbuE2bhc6kSuqYFIUUCxnk5j6zXuR
pinQFogh+zZGbN1AA7855ySxk84xn/cEegJuAV9Q9HJmb0kUh64F2sFzeL5Kq2ahL0Uik4ehFF+S
hLpBxOnGO1bzkf+BdJzfLoFP3+PzCiHAkAyNMJmSwB74C9KJElaX5Ro+p2H4Yv9AY2XJHGJsU3jG
XmUfjYBRHogDPBPBJJGA8jT9vUr9QTOPZEbqAGIGwB+nicuREpk31M4YJEa2wFrbwHZtR5TAuvq8
6zNHk8fnHWutxhODmjf+ZGpcceJV0HZjj00ElHf13+wC11iEGGFKBlJUesisISVkgqt3ZSo610WV
uAJ8xtOOLwsdKDQ+sF7L8DfSFmklK8Ey20ZqVzJwDStJtnE8Oq7tKTXL3M5GdSyJtY/4sNsmDHpu
xA2mj+MB7CVxI6zR+1fHsvXZxz3qkYGNpCHpMS5rLNUbe2A47+FA8pusipg5NBx/60aVPxP7OtKa
MJdPyoHYy1V35LhabF3Gt/pfvw7q1s1NQ4g/tYfxG/0ZpxX9vAy9sg0kXHHcf2/+axvhonAHVbDu
0mRehUH+CR0CrXOsoY4VrzEprwUE3Ty064CEQf/Csf1KUPOlj9xm1DbwHr1SKCtA4AlsiB0oQrFZ
FvqoBE+XIIGOkqD0VylQm4OzIYioY1zBEUev3HvYhUWnd0gUS++pP9YNQ7rg+a8iARMxN2dm4J/x
Yn1WMh5IoaP+Npbeeql9RuwdjEePRv6m+I3JuehMMmyI/2Yol45MJpXFsED4uPBe1rY3wU1MTHn0
Q+7Po509KePA2RN9tSameBH7W4M5uSJoq+85v/KY7GWY6B2qHLVm5590WkTuqVd3VXJi5Ot6Vfez
2CFosiNEQmdoeOzzYCW93et/4MOYDcP4kGH5d1MTDLE7Q1V6VIKlxe1eTE6RpUy+ax39WV+IDFPL
oQeoVpSC7KRIYAoQQ0DWF8NQckJ11p3Lv6eBjrnnUCWc0MAx1YWCap1qP0sVv/rsukTJmmrJZfiE
X2fWI9zYddkKqTeJi/dbqs8Jh9Yt1aZzHvJ4BmIdjXU0WRz4PbohFRm2qxRuMJX6zM73lXTbz0M2
gyBAjbTbuik16om2UHha7l8R2Rm8pvlscDWeOtNGeGW6QJ5lxRDAuuDZ5q+BJcGwEqLJEK6hN2k3
gg0Ul5bBU7b3jDSScsmTmNN78Dndfa0RjUJrc7wqZbJ3WxyGpyVrqRAc2sdciwSCb97fTEq3QEZS
1m5NpBLaVQx9jMmuB38UG9ZebQFpxl+0Ko1umP6WMWnTP4btYKWokezFaQye4KX543vF2vDQuIwJ
n+dgnPI2oQH/Ewr4LX4IHLBAKpcDHTCHkf50ozO34l2YKa905ak0Iu+sU36d+EI0fHQW9sj4/86F
5syhzhFBtGFLs03alXQ3XyMoopdDABjtAg4vL/4dct26GSA6JOlaeX1zK9hktl1cIbZ/1H4fdd6y
r20YlQZv5BJt4GOAgNOLJINVbjV7kiFWq081jrG9oxJUleCFhYOdmnfOJdk5bhXDjcZ1KFitkg7p
AVTLPgGKtQVxKdq1gE8BYHpmHuZ7UaOT3w5k+tzV8a5QWvRD9UiK4I9IuD0VD45TFX5ObCJat/cq
1naG/WkhgbQakw6b5AiSNFm727DXgkRBHZemhXmpgwMeYyQh1No+Mo4LQW3EghLAevlxOgSnoKS9
j4jQ1czYbo0myB7D1DztZ4yR5zx6/EC2UI8yPS4jM1LjO5m51MA0FG2EQohu9899v/jn1FhIzXRd
OOv+LwE27IUOqn5beBHN8RMt/WfQJ5j3JexKA3s5wHQDmLmJAC5rK6cI8axoqFA2Yu0sGkrRRMqN
fUTk0GM5MmGI1rZBuoAk2FurAmtO0159T+Guig4f2URnP5EBQ5DssFm0qN9G+j+xoHgxpSaZRCkA
AKL44nmuKfoBT6KAp1TRlwDXB2g3hJOZQuXxz48p2i3Cfc+RgeEwvM64YecvhiwpGe2DlMylhuxw
2i1n6uipIarjUcoEIJbDtgYobFol0Awgvsm3Yifd6s5WXqH8olS2Qk9iJ6vfp0iz5opM5nC/xwCt
cErsW8FP7dNw8vxFOwWibuZW4pPiJcK6ts9Mg0KjAIkn95z1b8bL7SIE8+v7VkHGA2HQUC+I5qYR
twBeZjG2IFpezE9rFeQ5TPjiKYloKuKipk9M2H0eb9Zkk9VZokmr031aj9NoBXaNkUNv8VSiFsfY
Pis4IBdrqkfC506SbJpqPA3R2mUtrM2G6xWrcsNQ+AN9C79y1jT7myBXEP1LrA+scNFHtbvOAzGp
r5Z3iJWNXlaDtwCLUWuZlGdeYH6mVxISj4gcLjaarwSrg86yLsUNQqNiHmk0WORO6/CcyBpBJVrw
gvcfF5ZQC50Ww5mptaUzXDD1KJfRap6iVTQD/XoweciX/eyQcvDVGKsFDtJKddK0PAIbNBekC3nG
6pVth6KID8HnANNfxjechiZ5utQY/xfm95AHTuL3ysat1U90LUk6UgH+QfhBsTb3ApXdBKJ2nRIc
gfZs1dwurtgaJs5r6qvkJ7p6y9VdjJeNSV37LQzvACnGCq9vFSBsFpHqOgUkyJ0u4cNaRJvVLTFs
vECTxd2nz60iueeilA4Kfo67LVQzrU5rjUH6aUHa10XK93AGXf1f205kEMNfCmoXe02lMu/BdUyN
n4MqdKIXnQ09pLlVSRDZtzVWFI6WH3hZbjJAtKxrbfyQv69+ht+HYCydk5OdDUWANEGOkfgZ/g57
J0zEs11sqphIqOGyezXF06fBjfEFcE+foV5Wtzx9z/XBx06HqtnsY3tl3ROWjC1h56C1vcuV/HRg
lW1ymMbIq9pMbqFwZ3f+/AuZ82Uc6LQUqB4sID1ApMibpnanu/8Afl8MrsjgCUEuXSXnAJCdOJrh
p9jewvwg6nju3hKWzEHk081GVhU83hnXyfojW01KTEEpwinBeaqPWVK/yel13SJuAA4PTvVmqmYH
umDW2xtWWa3sJ1tQOBVMBHerhE506XW7RVQeWOtM1z0ocFNny+iHVtXR41u7GMN49cLQIWPNaoZD
6MLRfsJDJyAn77GWjaIg/NvSS6Bgi1kM6KoyQ1tzGa4GwXGihN25hg7HxYggax2P3LjHlGcfl+Zg
UajIgORn87TeDuT40vSAyga83+ah7qpMnVOJv+Mis3gENA6qLihvEK9Tx/1GOkoh4Tkd885GI9Od
zIjrogA1aCrJlw0J435Y7SvD4SsDO6U6xatGsko03VB1vCZ4HQsjXftU+wlmaYOpEDSP8KJfOw75
XOTdb3SAFn8Irxo9dyx/yLc90WQ7rSE1QbcHqiWdLbvJdg1uVduzOiTahwOR4v4TQVket4gAfMKq
sxhpaVQDhBPHMLTTehu0ArCJaAm7fQDu9qtEM34uqV0hmtnW2ZMY6RqLSy6YEn9yEblHJSp+nZ94
fL9qewjHNVwAeR4OV/XT4qpfMtlrkef1nzL9kWW8S0V3JQcX+x3I1q2cVnYcxLna4rQ5w5CO6Hh+
B2wxB7totcMC0Fo4Q+VK7sH3UUmlRCWAj7EjFwngT8a82AFOsgDEFcFEGwrc1KKKs0R3hUvlYqbZ
CxWd4AL+3abNUN2k8mImWdHF2L3ojOHhAOjFydRO00GYz2b8IPKoUeV9DlFmLQXcboSRm3PWZa3o
5/GNJ9olYFrDr6WI5g+Z+1KidfWo07kwWIN/W3JoY7Yhmq0TFlWTUg1TrNqC9bMGpbK2pMoPOdnV
ENNFzMX8TrUCOEAKxemAzQnSWPqqrGl6H1pRpQkKzuB9M3fj7Gkl1QKb/ZcdhRPeIsYWK1DAQBGW
TR17Z8CfRPkuvUITQTvLoVIcQK+k7V7o4ytiex0ozi3vyDrNjs0Enk6F5dGbVMbjPJBA3YT3lmkc
vlnYHTlsHZLT7hFc5tYkD1fFVIXY3cT9t6Qx/Ccrweu3Yxm7Zh81eB9bI2sZukTRqgkAjq4Uf/Jq
T2evhew7E7dTd0UCFaWWQccC54g3NeWd1sZDMVb0IIumBCUj7jCOrBDiZMDk1dFfWFxOWyM2r7Xl
WDfxfbWDbHRhqkGQva89xl1dbTOuL+JjeVncHib0GavUgCpM2gt/TvW2PjFWNdgNwOhoxZXhfCFG
jrKqd37WdVWxaKGWBlNbgJC0jwHuiKgTjZGnrMxsJdCBOoNMZbVEJ3Evy5moNJnpMPt+YCDxX7aq
5lvJ790c4Yo557MTqPz+JzKIHJVceHhsJqiv68Xq2Juyauxjjq84QLh0SSPElR2PqxvWp+55B2nj
pybdsmy/agO/oXRC/sf2r0Rx/PsAs0/MgWKL2dDL1nJRG+uOXiENvswhIpL19pFvKz4DphQpqZPg
0k3thfmMAivLNy1bBP17HpzldqHqSLmJHzrTG1g4j5pDMccaIR2K81HBS47BrMHzUk8MDNv34Bqh
JNBKIXThWttkUBa0OCSyXc+9Xy4YpItbCBjSaY2mnCjUlpH4elxwH/0I2pB+mJztlVOPZWTiDfjF
WT2ODFVH+YWvgTaNSB2TNaWnuYrRq5la6WqgVYFAeBlq7wsNbEzzBTqddQVNSTkvTSZT22S7lKYc
Tawa1Ff1u2kYM4lw2gIrX/CjiR+bTiwjSu2ZDDjjee42YgCi8RMsVQbKvEi2pg96dg1FZhhFYTau
1TbmN5FqIH6W5WWtjq3OUg6fVCM/ujRRXWJ4mQtpXW07AGYhx+5mfi6PKPDKlvx66HY6FdGxk2X6
2IZwm9f8ic85QAskg3IxRV0DQo/UweY6ZjpkyF1dW3WB4DB/51Vcle3o9D2uKuQjRZZZdeFpyy7h
AUroVbr8v8acsrLxuQdIguJ+G4mySCjrEALnSSGVSBt2Q/7FyKUE5mk0HG3yBSo4XMDDgj7/Ck6n
ht1mjmEGZzJK7gKjaWK4rLhEgHhbSSoY4EvMwJ79o6hjzYzVCF535hyMf7DBXC0+Ib6DOz0LSygK
0l5JmH9cvyDYOuRHhmA4PLSQPhnSqZkdc3G7yzRU4nb5/0tG19xDZ092463HSRxottuJq3jaoG2p
rIIiz00ijTPPFmN7F+EwjbzYefsgR+yjDW5ju9Hf8z71tPIGB02vi8j3GBM9564icOunfYqo19CE
1OesIDyIuDQ5W8FDqIXH62U9ArxP0f/PZDtuCRl6FeaFZLBU3SlRjaR2XEOanh4ymZ4PlbeIF5WB
NAYSby2IyLEVbCDwDsbonZRXYKxpNo42KWqYvmw71/ANcKYLNUjWLkRJfzOJ5AznmUBkTQ9ImK0X
mc2KYJ39TSAvELgF+xftSWboPkOLOP3tt1z0sVjVhyN6YscuymKfLqHuvfcFW0EYnKHGRBTga2ie
NfqSVsbtKbE8tA9RjHoHk5fESpUH/fgrkP/XsdlC+mkEQGEr72RpyIyHiB77gMRsREG9IDMugO3l
2PjZEBpsq0QA0y6i7cUGITPNmdHJ5fe16Rklhug0Dc8zZpqNS9C6V0so7hWq+OLpU/Vo555zLnjx
3qp07yL8Zj9N+/A8gMn3cSv3zPaGeqX5ZDHh8UUuyHjWIeRd0oh6Lq4xXL7RXDCzimliRaLzp+cx
4ZDzEKtV0LGBxeyG8qkmPzAg3ZmiIb2fo2gGZORzVJAbhsfPb+JS8xyd1KX0L61fjkorwZs081jc
xzlnRsYMwaCRwtk+y5atBNHjyUoJPNrhhp7T0276O7fqkISPAmVVL0Uu4E1/f77T+XCWEyjNfn6k
7v9ez2/kFBMfxrZTBcaJEY4Rm2f89b8Iwt0wRXmLob565W3FtUIm+SsRXioTY7aPw+N1pMIG3G6S
YaW18B46tTiPFSYXARmoqDg9j8+8sGDV8d54O+OZ8DE6RqL31pJN2lN1D2tS9M3J53nL46u7obht
ac56U+2lAeYKC5YcgoFfvN4a+w5YXQ3qmeDZ297Y9mz/iqmJSRhN0jL2Biwr5vF6YKgZL6cXFWUT
/1GAZkRg6GRvVTG52wdV/27jYmzchRLC8t9MxIYmHb7ereMzOjIHxf0zs81JpRBOBgp1IKGRYa/I
dBGM3RkWPgXhRp676Vl6skrxFnvxfT4GxfBv+Y4MU7FFEqaQY0xTZoApT7eEhYRCu9ngEAZ6zGgP
86bHhgu+3d6e9Gb++ObfL2Q72fhBuxsJCAup0RU7I1O+AHUX/f685Lk/TCyk4eyCcPwzQb8FqYSv
PDtWKAJbZqjb5yPTjxufyngdDDFZ8A324GobiDF119l2WdNC/iT4A3igZC70+8QNI5i6lZS9iSgt
1hYLGLZT2uQdgZxTIWJKXVaimohFgEZsiOoNR3i03zX4ec7cT9e/qx1ByYwtUPWxUgAgQnQGMnv8
X9Y+ne1aeWKYSZbddZErloGbuOweQd32h7wT+bzqxUwOyZ1vUiN3xfSR+7baEeCaZ+n82NoLdBzj
11WnDlK+r6keuw6O83cCSU0BCWdBsuzVZRcU8C9gARDpcYVJ8SrGRyHOjMt7bjvF7SNqg+0aikUh
L6HARSdyvUQrqg7x80xP4x0TR4jhrHjfJf7N7dnpm3vx0X9amwdCy5tdGIMd+DCKIvsVaavh/DVG
uV/i+meedVfmgeSRrdF/dZPVZDvs8CDWB+gwH/LcGWRmJfYjRQQYPLM9o3YfLgmtRZCIWijvLZog
R+K34wC//Z31HCbxOAKk+G+6S+I0wa9bAZTTB3StKK/nxt3KDrLAE/uGbPKDayKdOIbunDYAJIjg
czJK9eTY7ktmA8QZeulCtAmob3hQkf5khZbBEiNU5Coo3PY20fpZ/dFlMeEsdYtaz0SAvh92mIrS
6mjFGyeDQ53rW+yr1aK5KUeuwXRGg/ozIvPX85kC3H8VY52btqCVHtt7A8f2NZ5Wm2o8xpCQzVLX
SLWSCVXoZtQzDxQwwZvaXFCmBOCRTs72cn+8A2MwfKt1Q1sV/UjFjGR08nyYmxNmOv9GnNL20Mdf
HqUoI4fxM0e9TcoiiwwtTTxKyQYmBDTLb1q25X4n7L8v045Q10/chaCXSz1gvaV9034EN4kp+ejb
k5heuDBaWwhmJpfWL//X3SH8qo8RvK4W3YhwPeJxcb6838geWR/JD3yitDSeXI5nysL0sLfcY8TI
NKMYTDIQ7qxHoN63DuYTzvbQg35iEeShNN/iN6xjEGd0HYv2NHPtIiiiPcroZTyXXm+Ftl9zMjxe
tsYeP6ySK7GSwZpbqBuNioQsBj13nJ+Ox2Iw1QdkGMYrijV7OD9Kt9VZL0YesXnfsH7QAPkwDPe9
iDCL38Ks8GuajDnkQWAOhPfaZYTvHWaLPq6gZwZiyKXEEPIdy70r3Wco5Pa06Tg124QtWBwsa5/t
JZldZ/t8qYzL6IrDTfhgPHrUm0VIEsg0cwO09wpBhfs9UxALIDIx84f9wb0dx6sRMLkDT8Yut5cV
D2NqVw3FOzdFaTBTOhENpY1oB8n6GY+7r4Lcx8I/uOTB5sJeODVzq/absL2heYxziTXnJJBgssbR
oFc/hVOE3m8cPSE0vr2eVCMaSzB+03K2cy76yaWXcsFa4ibwCiWHg3RuIltBPdf06b3paPuCFsuX
OaTeVniD2EFF4R+QWvQwSu0PgJFmNa/UMB4hxOiNZttyJJcsM2Bhg5eUDNiAhffaoQ7v2XAl2WO+
QlpOpI0TAxPTS0YjM7DcjPGILABypVLnnxWAfWpEthzPRlVbq1HkwIk1sE0ymmIq8tqkdQKdPLtF
3B258W7MmR1JL4WczOLcXuvJLrMepcNMOb/GrpNBqPwbr6L2oXZSjfVfqGYeaZb5ApdHydHBy62l
WMQAh/IrGEihSZfVlmh2um+pbYGytn5eJ2petzT6loFR5utOJNSgIUrFT2OBHErY0MyrSFtfV7bK
p0Fw5b3z8VWqrD6HnRMLsfjKwJIoRwSKixm82d9rsLlfClQbAQivTLl/li9upYfRQmM4w/G0ZNEU
kWh53OsKAfNljIFYMQLZ1nmaWNeYP3UbWTEQWEnDr8MXctYZnagN+iZ1RNOX/8X3ttUkANx1/GXk
oI97Ydgaln3w/Rcnmy5Gh1v0Pb8MKZwqGnshLokrBjxKdIMxS9ZuCEqOjK5kAlB/J5CX9BN+UUZp
54Ide5YTjsa3zJilQFHGU0XdOSLGyP5jHCYQhMsKTgPuEij7K3v+0BYLcKViQil+oaqOaVSclt6y
IICLqXEO6D3L6VwG2IFHwrbNy5zGqF0asYKKSpSzByM7Wm1THPQdWJGNUytFPFk7sbntrlich+Sk
awhEPa+c97ggqkr7/WqJB/Q3fku1160MDK84QRNMSta+3v5CcCx/XEtbYkQ2EOa4HoYWz8gCQ4fA
2bZvzeLMgqlSDlBNziKF8pgD0JghYSI9MkKcoSM5zHPpSdgeoDL2DUHiIcsQdNBY1yfqB9UGpIRf
E8hdyGRnm2UOr5JB0LTyKhZU/McqpsRaj9v3IpGPYfmSIqyzPIl5QW73PDQtyq+iVPephfeRVKBR
QowZo6QGxXBVUILzaAyOyrLWO5jrCvCpaIiNvaNFlsYPVuhgb4JtdEpf9pe3Jzuv13LoK52osTUM
HA9p8gJk1uneuR8xM9H8vFl0Pzb8C0xSWeSmnRaEDwli7+GMeiRkk1bbpMgU4YW0cFQnJVOVaUV2
BGuIYYons6mqWPKGRbNI8t+zwSpzsKHR0c/wwp7KKkuRMIijF7iAdK2Z1krfcTjaqpZEvLlBqmrC
uVGPyF00bI/6N8G2kwZr50ivzE7Izw1FotXZUFeni42VIZnZC7xGF+qGXAGzxNTPAfreuepxC82x
0yBXUKbaHGlFj5SmXuSR3MyqdXdybLfjwXhXJN6vj00E2m8cY72K3qaoOH2PEm3NP118gQJ2WCMy
0JQIMXeq3D7b2fTkFrLQjbMItI2DWzOX+bgtJYgXAPBnkBDnAy4hli8oNtn0+n71oRkmQ/BFcG9d
Br9osvZTwBrtPSnOSZSOE0xQnXkgeHHXwc9NPznsrH3XenoQ43qIzuWjP+HubOg9HrO+XRgUUpZI
ksfw/wbk63OnMixQ+JkHpVnFdu4cbQb/QucdPvwUBeCMNkIXvDEvzot+ys1HjuE8MwUSBf0y2yjJ
w9eW3TSpyEeuvqrtoK9fxqOqa1YLvvbJZfI2n5OvRmskMgTzhK4qoqAYxPzhsgaKFk10I3f9TMt7
Z2iOtKlG99aM5keWNbw7sb4VfUvUQo0BI3TbIBe7RAsh/0RktKo/3j3+HdgG7cns1VqDkXlfDr2O
5AK+v9eW/UBqruOLJqYm1pcrrZdYDcM2sCeFO86gRzVoPeQhLV3A9N9T8oiz6iP09ij57yisQueD
m2c4gmctM0/PLlcBzVxumJLW92ah5jnXGBzIp4IIpJQ3oDARgKfMCqnt2lj3+TMJoNcQ4yRDqHr6
g2Jp2/o/8gEIaaUiGV7eck/w+oDVF2dMXi6+fa9M6xFQMdCoK8sqmfwvZAU8ICs6h0Die7FgcxtP
j6KrEeDwZmmnEdOds0Ae8uNvEAu+A9ugvxxyzHe1WUGRB+/uwyMFxuvQGjno1M2t8g1D6j6EpFRk
vzYCXSjxV852BjqI7ML60HR+SElck24713ryyYFeAjUsfCwq9NCruaUfxWjy5QWq68FWWAteA3so
vIgUS0kxzrnnAUYmvvw5ymp9GcKLIqctRULkN7PldV5l4LgymgD3cD018FZmXaMIqGIc4ZsN6xbn
GrYaxyYVtM7CjVeMMI8j6MWlIQf2oOHELqT4vDdFeO6NUX5CpztpcJZ3hcOxaIkg2R6j93hLuW+q
ovq5PbwKyh/CIetWSq89WawJ4s/nd14gGLqPfwq+hXnHFBB75CalRZ6UIyVUEIvyi8QoWMT2sVbx
g6Fqa+ofGFjHkrKFuzT0idhutnoF5aSvdDACuDfl7c8ToBb1Q/KPsa7iKaC1WWFbGeQH7o2jmwTM
RfnH8NFeBEhr11QhoXgZ9kJrZbHoXI6fNNhXV5LCLlCtdaIGxqTrP80brsXiIpoZljUk5oiKxUoP
SbvStzQqsBvktBLAaLjFOK3SAj73umE4IRewUxVuKnpE4QiFIgEto751g+ufMW5cYvgy4ARySim8
O/g8e8EaCHYBm4JYxvBXcWk+QrlXL91ohzqePViDYvbvN7UP5lGAIKDNJOTtc7iBMRkVQfTpFiDL
Kn92htrGoQbA1Cd3hoF97fbzCf4I6CgwzG3dYQOV838kpvNuUgHW572dIqIiJCyxtNKIT/sbKq20
JLte6XenqaSD+kaG+pi5+eFbqa958I+aNrNoMhH7KzmcYh0pWpCCld6mis5xnq1e2u5Yk3O3JcEl
c25iNjih91B/6FjfdTFfUWCkyc/dll2HyzITWHkf0ZVIckXlh29wn2D549p0HZrtXyWZ065ByUB+
BQeJeJI8jHUAMslvZz5ApFv4GselbWi1xl8VwBbw+NuUqhP1kXdrQakqHB9/TjeA0uZgVFA5Rcj4
b8s2gPiiAOf+iIIMYSQUaJFhYzpn8XBFs3H8T1+TQBGzDfhfaLejA6c0lwforCNX2/Ti1jbRTLoh
TZAYy8091WUlH/sDt49bxeVyaENljgGnhSxAThEPHncMmoMSdfgb3djg8RI6QNlTzW9q1MCMAI0D
tDSsPJpgNdFroebHfMR8+AWhNi6p6/TRTTL6H6ZbE7GU46Y1rkLA4gLObV5VI1+a4d9HMrEOg9F1
ci2pwNRjijSqyU7rg85xXJweqt9BRJUAdJn/4BpcdJqg4JVNK/Gk1axwjKAxYxbGwpJFoP2tzYph
42+ebEELup05pR8Avx1pNMA3VmkiCLr+SXkJtzlpWc75Q57oG+ajSMEEXRtXzQGCa31zELPZmxLi
1Yhwe/f22yMNcauX3PaOC8n+AcmLsWKP0vqwJC90CU/XXf4eURNkqQcQf79RjXKCRyKBLoOjD7a5
aA3+f7VAKZQEbW9r/hGyfQ+Nocn8MhMoVA/8jRS6uYIXof5Yj3HpNt1Pdc45Ol9k/j+RmFLS0zAH
RRkFEaxTUXChLPhc57cjdDYCWC51GWMLJr/uCCbJi6BJQlVd39PNG/ibDWgXr9bmBWCZTFX2ZByP
dQRW19V4/kb1YrxLXHemxXzWHCUVAlDIB9GNvz29ht2Wme5T09eevBPWptnqW9082ly1Eb/VEECU
dHGcBRM2lxJsL70p6RIXVDkdNHyq+xa2Rbtmn/goHCK0qQ/qCP85J0v0dsaeszUXZIDTnLWczgiY
AfbcbGYcH3t3HPTM7nTxbLo+/2Y39aofGrTB3CcOy6xsb4lZP8T+eM1Rued2MUlfTrAqRNZmC81g
rZqsfKe6hw3k6HQDdOG18t7mrPtg2SRSyrYVvFO2oUBhPq02SNfiMEJkabr/lEkmqyFHsq9VFLGn
QtEtqGgNI5eaVyeqRpb8defiPLIpBGI0xs9AQcXjDHPdaprUiVzuZtIAiWsuVEzyomE6H60gKC1P
Pa2rjcXGmivV1UskFeB63OFE1myPsc5kg12ONylhVosLwVCo4ZyXVRgMih6rmVqvzxxZZ8jTfVHx
nyolcbUcFQ753ywQ9r5GTqE0qxbNnRJAF3h1Dr2VFf0dA+/xdDhVYRerYJ6HvAR1CciX6OESCMGp
IWPB0I09zyvzpJJE21WupqQdPtZFXjOo+59eAhN2oqPeUtnuELq+vaV/xVoZkv1WdfrEDFLn+KkL
MWeXc3iuYeANOOe8JwGOvhPqTpYLrOW8RluJBBvDy9HyMzvgC0H9u5xfpNd5mrxmFdbmvvLpECiB
l3An3/Xu8rX+hr8HZSXucJLM9rtteHPj2OUpXzHOD3BK0/EpVb88qNctKFHblUp6M2rggfj9sNxh
Nd65+S1okP44QF7OnfiLxSQwrp+eePXPQOMw/VgRGXUYyP+S7EoNjl/kmmthCsPqbGVXFxmdJcss
kasLLbm6uGnfwzB2ltGlGmlam3WOwCle3jUZL5PJ1aWygzvq+9uuXmmOgc7t4cOyXDMZzWhwDN+T
hONuBxayPzqI1QAtcHEFZZRkHCuKwDOWoiSvWxmkeK0uvrIm9sgAcmbeNi3uoQWMatw6ig+5X4ig
kuahML/UALTIOoHizLK40+1lzZpOVerOypHd9zpIrro6L6bsT5pdw4okBIbqu3zcWDPXuuEOi6nf
SsUTJrmDkmN57WaSUAtWuQPMmt7CpNT0ywWLxnYUPtFhXOu8QYvP3mG8E/0p3xs7zk3/2K8WP9nW
2BImmn4vR3HcsWLp/3CF825Aero3cTl1P6lvnlpncxc5uPJjmEaJrdzRrnS18GjDGOfBksAzDCD5
8gZXoP0KiZ2XnHQFKOIug/imX0plVgy9LS3WtQNf8lKvNW6J27Q/uUyoB0PDC1IEMOTdOtYCfVUm
O6lq8eIr0LGdXuQByHPAtMZyNF8X6RDBS2FR0KqDH/qjFGd1/gFpS4xuzvp66OkMrtUTJW4YIzFv
XOv4u1JjjpJ1xbOBAYzWJC1ImLV6YXkEaSd7ZDbYn9tkDXQ3xerGT+ZrGYUkSChMfz1eAGFfO1MS
NmVYX3CyJ8BSIVoJr6CIfAcjfQ2hYn9rmbBQl8h2eurxPNEJbHiBXS4D7TFb7UjEROPyijGd4Lss
lCtTOrvF8Id02wzfS1b/MWPP9o1vr5P9KAxevOayfLjy8KmrgKupN48EOVWxjVxqHDsg8LsYLzhF
1PQgCaNBlC2ioYDjGESnXCeutviRGtC8v5OIrgFus4IY3TnIDKs73TtFUlnXp58a2USuGknPjf5G
p9pQkMoRRvPMFsxYH4pGfKNfw6wthjLNRFEPCPCUNWJAVdXR2ouA7aAw3x+vs+k9f3vsi6i+aTzK
e+0240MYjHNyqJKaWJxmTxotB9PXehxXiZLaKqWlg8CTVnnax911zlNBOHBcYSJkmKh+8Jaici/h
AjIUVgTJGyqsxzH23YqUWuXUPL81ZaQWvhpNJRw690W5DunJ7fF/s3YWHti7hoKWLQL870rJQipV
oRgd7Kvo61t4VK8DE1+yxz9lqIP7+Dj9nTmENOw4RfS91ALa4lu5nyPuXIHV81kOemlVexY+zyEj
m6wWcxvoXuhZGEFWHKFIc6FAaE4xdpd2A3YKzNfMYLBLXw6aTm2PJcjp/xvj/c7SNRqozqFv0I0i
oZZ1mzGQC7De1XOiVjpGk0F8IA0db2G2LZDf31ule51MGOM84k0pqmjTWp2glKO0LKDIFyc1V0Vg
2AMkaJCE7JvSvtjleep38zKj6zq2MEpP3pBIuIVSGr77sd4yDhUuhbK4SEwSE5+yGmg8u14q9+Y7
z3UEwApVHc+0pNJX9at0Q2rlms9frUEdgiP806j5l4Edp32vMj1SIMF0JT5k+acHVwrw8E/o0lAA
IsT9DS5UlTpmi25JIf5TKT38hz/e0TGUWqtpO4f0pFhvqhVEz/F3aO1kJOI1iU9EYbJ5rM1auKIp
XItogWsW+X4Bb8UEzdf9iS8V8sQn7l8GWhYLIDjLpQSI7SsFXu684YI07Cb977tjXh1UCXc/cgnl
cA4jbb1uzG9EwBgYoOqCQ32wrMeQby1fEBxqztz1OYT46kFzSuEEZ8dlt/jpVFEcHQkQpNmeyORW
kDZvZF8AeEn7NzrGG4mZY4b7ScLZX4wvBMH2AHH62qFTx6WMW7tRTGkIWb+hnONxup6ROXO6BZTT
6nzhYMtzYjy9gRJutZaCbs6lJB8p+UYSMGRbxyQnNHrb1ZrFzmicY1a6L+co9Q0Db3pesibexCah
rBg5RNkMRl6wMAJBqFMrv81qehffDzdm8dW588I8XxDGOqoGNtKqxNNWobinwk5QwivfDzomg2/r
HJEl2QAcIFnOPzAwkQY6892A1hRz01ElH2NHyRX7UKhu86j2e2OUFTdfnR5NbXYxVI9g3Y6+O0Wp
NAoZebZ42fq0aLbKWGly0Qh0/ZYeDRmSHDuwtCL+DK9uMt7ojWAyUFINa0DgGiG39Hsf3OGzcWey
8Z7me238cXx0GlyCF6eQZBsow1lr+SCGNJdauHRgrA/Hq9Zprr4Fkn0voMBprEiWO1VGMA5aTW7u
gIpUxxmh/SgJfmx27xkYYodGDorHRFdYOMd66bt4+xXJc7pgReNzSAfCr4zKetf7RpmN+3o2Dbfh
dxDg4mYbN+gIOTKOPYWdb8jijn3L37Maq1akHeCZ2ACQMglWmsL6KDxVOI2rQJLKGeulMUPX2tIN
EI583HTg+vhax1KTr4Frfnv+tl/OVTGzm2q9x9LO3oYxKnyVZxxT7OqvRwwSGKn5fMMqnTtyF4Uu
EE5BsZRb7kmf7u8CODyeg4GiAzM0lUpBexREBt3eD4XftP/pQOFe9WVbIPKAq5+zskZ2tEFZZBFN
A+a/Sywz1yTyI0as5Svncqaa+iiw25oMNwjaAR0OkHc3s4unmYqCJonSUMm5VuxKqHKmULVTs4ku
fwginFjQg8UM+YOzQ80E5uTa0b/SGI6nGGE0Z8AyObuYqZ74+WXx1U7EWCwb9P333U5mvTmMmsPh
w2pvpcHJlr8LAexZCWCQa2GmKPfmoTUhftjFP8PWjPwhqUCutKsmWDkARMnewx9mifbzz0nCqRdq
vZwtrW7I3J0P79QorU0s+N6sq/wJx5pqJ1KJlN1Rzq1A/a4Jr8KB4W/6dPCSeWTiwWuNQwBR7VR2
p9s9lsunliPSJtXekz+da3BikkzpMKwdjAT+JV50snVMNyS+Re7IKziMb8iaSBUGDaUGncOi+w+b
LQiRZ8i1PBdVD/jXbO2LMNXa/3KUB7fwopqb9KDT4XTt49nF4IuWRI/oae1O1BaSSWhMtUUOLNEV
eSqx6aq21aP1MMwTI9MlPWYSz3V4vUsKI1yjEByWmrnJFM5+jlmDgOmpSeCctM1YeKzK3n3x155Y
bNuTaxAOCo/KHghWzs5WlpgzbMqf1w91Ds7uohP18MYLhZp1BP9yFLQda+b2pBP8jBuTZ9btMc6S
SYQfYQaWxQn8L/bnnowZcZ03vJqEdKF7cmeGPUOX/+e4rDFPfgI+lVRt1IQ6N9zAzu0La1m5T/Xk
hibvpTL0YOPK2weNhSC3SD9yV/NZLBwqQBoPZxdxxX+dhQFEQK1OrgGsB1Nu3HnsFAWQXrJhEYj8
OKnvdzNfv35mphJb0TrnPawz+2B12kh9VDb0UL4N9fIYsyWy8Yb8Un1tvjbJDa90M6cPaxXuHIrJ
iRLtUPEz9YRaOWGfaZKIeplm67jnCIBHtzqWhB41+TGHo/kkwanZr0KDTc+jbhRH5BAHp8fCocG0
fA4C71SVxYWQq9RYiEvpfb4Hh6SvZslg83ygF9ZOgnTgwLWQZ5Ouaq45ROSc8s174bzbyysLERSl
/z48E0mfdqhcfze+CkvoDuNVbFfiKdSGo6lNZ3KyoyI+mRPlykZ5rJNyyQVOLQYXnhLIOgtV1T9N
Fuu8fjgzrBfTk89SZVJ4Zx3JS7xJ1aUUR8hkKWnbhLlIYTCWUryYIvdf4gX19e/ukUghdAX78riP
8ogYhnK7xT2gptPjuzxylr0ehS25qL4izUodC+8l2QWJDA9/O1+ONXn7qQ+6vtCWGHlf/jcsukIB
ljEH4X9ABFfySo+1uvH3n4BQS1BXNntihYFlxQdjyYM9XdgMZZ5Fqe04CjQzh9QoRWQ9OOHHNslY
6EusJCgo7c+EKEvMMHB8zhrV+px3kmeeCODp5ibTiZNykCdlsxxMcTTHZlYjiX1/UEYPb7AyfSNf
7+xYb/IR6yWJhSju7Sh8Q7IH6F4TTsEDXp3oHn8dZ6mDLjSHgVBNJwg7dnDQ70//SflCcBl+yRL6
lQ+CIfem7zWaCSgTe0uRGDcmpqKQH8N5grWJMGuCAPMypYPoYbzi7G9gyIkzOrym4uYu4RRk9mNh
kDUMogjp39mdI0759nXpE1B1HRDiR3y1B7B2VM/S2M6r+pKskGuVqP7CP79iBkXHApx1A9TiumN2
dMT5DgWRQhoFcjWBXn7FZsMsYN2XJTsUHcChKJxsiOAWJzVglTLU5xIAa/SjH/Ied1Yhkn4k9MGQ
9VCWADq2T8a9UF4KxzcV9GpPZH1H0L8HXHZ8H36jV2Pzsgody4IKM/bL13TPXpaadCxD5i0Cd086
1YKcI+fEoxtncxWTLuP1n/u27gMDmXLMc4X1I22rW7UWpzKAssXSN4OQjd9jry8NYkgcs6vC+0Tq
GOhspILtCU1PRv9Esp5Xn+/+Q68FIySrqYucM252Jf5rAdAyB1EOPgXiqKUJZRs1uMGbW908iv9K
mry2RQjobnT3F82a6xGIzCBAw9mdPZkRbTepjaSV07rzB0WWa/0ipeHgz0hLazBo8rKz/RXOFdkq
+AIjSHWblnMdn/unkCTAHKIdECudSoOdnfmTrx+PMES7SNzZp0Cna1xEgtdONNZbs23Di8dOe98u
FDxU6QS7K0Cz/YGYsiL7S2ZbVIRJbQ3yd4OFRksnOmKQgYIdq8E8ztYe9KutNF5/lhcNQeE0L6Jf
QmYSde4NeglP9XdetEMK7xXovvbXkqb/5F1HKIIgw/bgoFlbd5JPcuqKx3YhEcLil6OV2G2GwX9+
0tmF1ypKCCwOKF4AlEURspKTXTqDkBkKaHdInUZ4vpvo8fLnh8ZR5eaYKCrNWn1i4YanQoOtDyKt
UAJ/jz8Rh0BazTRhbdcFZsJad3Pg+1eQKSPqAu9aL38hvn8Yh+JR9Qeq2Hb3y36njeqa8ewi/TWv
37AQV6lIrW5lLB1L/O6SLnC3MRc81NoHIWf+XEGuTGSmIW3mRj0eKiTJs8cjewQgiuZu7YZxe3Ks
RV2jQA89q6sy0zcA6pZGmKdAtX6F7gZhbtzBOZeTZp+DGYywkw6LfdRW4jWwEjC0UmJ+Lvcz64Yt
D6ul33QijlBpoaU3TG2oex6x84cdUT/efCZStyqGK+75+VrDE8IGoaxWbz8sxauumpBhnWcszhOg
jTIBkv9UFBYi/aMq6JS6ySKZRRXD/2uwTBeWIEdWqCLvLdnC1qGG4yVfy/nyXisRMiF7YGQZBMud
hhdFx1rfIF3Bb66Qql0bONZf8wsCmHQHIsgLribF3VPpuhN4IIhhLws+2sbnApuOZgNwJHioqea6
v6ukMpyy5/vepZh8W/wSZ35+rcjXIRZ31t5BiSSTiSSEFvpywkP4z1PcqUcAnVYjd/numtS0bBU5
4FIXK+SLcg7C6AufMJYEEBwVSJCl8fFtqfJINvTDX69ugWqMSP+eaeTsJiNB0CMN4TrVRNSozYIg
2ugMGJZBYAbZOOYAdHMexAO/QqZT3c4dBOQpanmjQSxUeyc0HBCM97rdXU+AY9sejWN4YiywI9Ka
jUWt8hQ3b1VRRGNjoTWu/L9fxu3Sj00CyzafrYZ89eUGm58N5iIFRYFhN76lXAYPblebmv0gyVld
Rk7+iIC1AJNCdg9HqbTdTAIjUbHNpjrn0Gb+2517fLmMHIz4VyNKA9UW2ZllGakSXTTmfeWbSOB1
vF/qnoYZ+c5aTsaUZezb1A7S6x3soF5FQA03BzB1AuseDNcZ8r43Z+FUI0MrJsrp7nUkJ1ONiN4M
R77vLxCjbXG2E2CHBOO/CeS7uZmksyE4ZsWshgRFt7W74EhPWXsOwe/xuCHNjAs9JDkzX0egOX3x
U1HTm46O3oBvwDdLJuGSdoiZxJuUE0xkGjELvXLrsAmZKn6PHodv+XQZI+tqo6GpKNLAuFFbb+85
BsmBRXUeuFUneEGyRMGl2ew62idl2QtmBo7IxLcLSNuqMbVY7jwCX86vKQD62o+g0tYIFVXt7bGS
gkEBaj39LJm+IT671dANKG01wbfUyjhCMBd0X/QpYjREAJFg5Z/f41riovyM76WWh9lDdHlKjJgE
/iwUnlWKB9SlC6TiBq5gpLqHuH7Wyu7w3tAzDJR7HkQEjkRKrGJhp+pPngPTAT9Wkb+mqXahlSp7
Kpos42oFhta0FgyZPZOsP4onWK/51MPH/f6CX6dK9XuQV3ttih88cD0MoxOEv70YIrCJAWK6WnwJ
Z8E6Wsrouob16B7js6J9OJ4wJkB57owSaRBUGwAL82L1Sp8XfvRmTfD8sC6ncZizhhfaxbAn8yjn
787l2NZhjBznq+Q4It9p8f65rO4XPAPdNpdaVy7lZ40MfsIsz9dmpLM1RH9GFbqhVbWokMurOyuP
HQxI1XU/odztj7+tIZ7nMuRwqFI8K4M5gRi2g/U4mRx18RFYGsec09b9mn0n9BnUUGSuom3sn8K1
Bed5/Cc2Byr0h/miM66UdlD5kEQHSkxzN8XWvJhAyIsn/PKk1TMJIkgOHpYtITQaGawfoKZLJtaL
RckZINJXNiJlz096yRDLqsOQgKluSFVeumb3VkzICONFzVY3tpqHV0o3vXJxCc0mUE1CooF+XZAp
YSlWZW5+4E3URhGbXtfxQ0xvWvWiH4jwSUBELNO2HN80uI7RNr8Ca91dcRQjt/3lzOD57h+hB4VX
Ty2+xkgRNtwqqNWlW5m0csK0puQgXrZ9E+gC2aHhu68956HlZ8u2881qOwfKQxaIDipuC0BN2fpo
JoxMAAss9WkMBSEWc/lQX8vzvDCutbpJjF32eeUC7tnGwU3gMtMlhjgnwOJc2LfTATNJcM455QTc
kb1tUXnwTAkbTDlsWaD6Hhu4wtugnvM45mpyg0yttq/iCctNzA9QYE1/tB4RuxO10UCZtoOrmytx
bxaAEqS8fiDPy9LjT6cjAoqPogQQ5Xb3DJICh9KIM0niZx4y4PD6Yga+61Je/ELUqgjnMaT3HkWU
GhXnfbEedJ5yHUlMXh+dE5Fo0L9JXlslEgvH3KWMD7fHXUIUtKjEs+Hhah+TrL8O3LePsoR7xlFp
lh7b64rF2e3f0A1APFgMjzfXiOd4n33lRAp58I7QF4j4dDNQHN/r2yB9Vu0IRDK1CKjQXZ1ergnl
U5UfVuhmNjrSP6GhtyKKbw1FTvqZJLaS4ptOfVAcvGInP6ht1q2vclvUCe5MhJgUCzDkqAAL6+sP
dLESMSUsumIRAzfyfJYtis4p5EC41c5xfsDoSt4VBm80E4oSqRoiFMWfloPGJkWi2WyrrSlqJxVT
A4MrY0K/WMI17plz3iozuFp1txqtRsJcpz6o58a+abexLbn9n/1W0fWgagNkhcxki2iQ6fIhYjoH
IGrfk+DgW6v5pI6elMzsIXRUFNSqUFdWPdP11FkvOUR4qcImI3pTtrDF6y62Yr45PyeKA0iZ0E5+
AovmWnUzTrTn4ZNX6jH34KkSrrum8G86Z3dsekghWbTEevX2g18miDWo0vJIEL6M458/vSnS2Rw3
px8i0jsBEJUzBqxN30ULmfYwQSjBNzohjv3lLiExop3KSZJQxTQmNzQN9qDOmwqCKiSf7p4UVMMR
5gkn+SGnYqVA3L5aHL4mcn1OP8qf7kX2D9AbjYaztn1PMzFuTbtE+QVuPWyw0JsmiJmT+dICK9z0
sVc42ouQl2CGtXT4rBu0uaQESObV1mkJIOVkwyuJwO1XCBMM6tWEWm1HrNV5ofYDmL/zr4recfid
1Gv7MXu58+Rc3Via6sbE8merZI9PbuItajsXCTzWEYJDzEtIGZwVzbKfiM5tyfLpIOLg9gIdGzLu
Dl1Vcg8Ux2YAVOjtQ++Wsmf7I14cou9aU1RHZC6wqUGH+j8H5ri3GjzDETIMQUsAZtd+VYiqgqdi
TA96m8vewODL9i/UUDp8Glvd58AKELhkeo/+owSZ/YObUfZ/MHzRKH8plvyjXuN27BYevljBDArc
6fNs07kWF90WPioM6FiFzc9yoIw0zWAedWdmSYEv9wFATxVePm/jVYiPYcROUdEkHKHMq/mytH4U
4UjV1kpVdXxC/9UW5G+i0blg//QAa6E57BpQG3FcSqfJaJ8P9nMQpmHbgyQAwOqakjoDLb1Q9Mx7
ZraXzGkyff81cHxY8Kw6fgWMctGynA3UfkH+5CtYA6kyNJ9VqSmRSRk8+d7BzUHrJsxS4KMeBZkS
4Osm21P1opl+lsfzgZPrQe6pInCXIOo1recvMpxRmzxU+YYrPMQCrsFa9o3B4b/tjhjegHXv9tme
dX3nO1saTJaBCetZ0P6nCNZaDXC9MDjnzX/ekbK+CGoFfLxYN1v64BzOkzx9Plm/N4WNttxeHwBN
+5+nCPbkZVQROPLPflNqzftDU1thE0kuhAdG4WxBE9HsD21sIFT3vJsFS1Ph0/L8QGE/3Hh4cAX5
YBAP8zJEoNPdUGOLhbb6Ig1mb1iBmYiEgFCppySx6VxiaPRCLQer/vlM0iB68BPngNcEbL2h5aVp
Logpg8sBZdHOsYXJOhU64q5kFPI+VdQWcOhkilFwJlKlAPjP9fj/eLEHpVHO64b4e8bkvwSFy+I7
3UgmgoH0+faL1e3elzr4WbPvw4iRqca6iqYrEtbeBv1h7tcfznA/7hH8595ADOYqZKWNcUdeW5eA
wpE4V/V6q5WJjbRrXLXMWxZebpif0e4vKrJAkqS3TLxXjpX2NInB5+s7hqp+gzCjpVS5b4W0Vkch
a+q6sQjYhT2adWHDql3KADsae1zw0nvKLDsVN6laVnhGTsAPDAJxYDJ55HG+EwC0MjBokosfhI3u
tOEZeAz8Ey/k4qOHhKSHBVOPk8BAfbC5ogGIZkyJhvKGaHj8Wccc+bb/cY5Y8HkdnjRrTOBP/+wr
qrDpcXq3QVYV0yJEr96PF2uKMP//5F/BdjiWMDsGIEbm/dkxv/cCJEeOCtg9CcCcPNGHSLaqt1jn
uXicje4Tgp3gj0Rg7Va5StvWjSZ7B8+FDwSThORhspuBu1pCcSMfZrY7j6KyGUeUcbenwoYd/jYj
jMPCiV4VoCsm3qmiEw1PhwvfQcR66GneraZffly+VBlMPzx0Jc82dN2ooyGxB+gsJunLBuVr643x
hf228UD/FvxtCVux9oY1U1uUTN1VwKT4Kkw0riYwNhYWC+ZkJr1xeUat9tlW1gjqSo590L6AT/Tw
Jnb5fBYJKrOP2IVyxPbaLszPiZG9iPXwJzFYTtmR6Gvesrt9M3gtN9WoVIN3A+Tjk3PCVaxWsXxY
xeKjgB/k/UqSC0OffPDV6rndSaMtF6YfuDkKRVIHxvY112uTJslSUzpF06qq9qeLKYN7yWjy9CW6
0o3cL75va1GVBj/tF1wN721pXt1IK7pPRtn+ax1O+YbvKpg8IUn/fpYh7uRjocRw9/usE/yKhbUj
PfXgiH10segvTCQaC4gyKDwgIHTzXIZVaYwyiSEooo0yr9p5snxCWukYQlEOv2yp/Bqr5n+rLWfb
e7zIqyWedNFaSbLU8m1SZF4DLbMnxH2/Qev9PNtAEB98BgjAP/zMilRbk2ZrNfuhzpu8dua2D6C3
VHwVFx7qM8YIze1s5LyZsbs/BtjRu38UXo+UEQ/vNDhsvs2DxpXJ2iZ8gd5IysprQ3Okt2xMXEk8
MrP7qfONjVoCgwGXF9FFE022VodbqeS+dtQL3ayf36FAdXx+kllSsR2qBU9S6towVhLTtxvbDNLP
joG5bCwmtw+oOYMJA3l34xPzETa/J9ZQAeyC8Ioodt4CUtOvJF5kM/0i0NbLL+SEYbx2m25UjT6C
nnayKrQW096dqo7OBuvRD6bUG52DO4iBdfxEgQrHjyQMHANYaQ5LZVWgNn/umCPXz+ATz0p7Fus4
sDM1lecFnA1ZQmfNRJstcxu8msfelZtBtHJbZA10XECmSwoQeoKtW7zjhYuoxi63mH9kTtDPH+UU
BpAPUzHaUhsn+Vn0DsLLXnl/pWWJGSt+31vwtTdb86S9Mhiq4NQQwgX5vI2gUAuHO7DN6O71eM17
gifhhWG9fqz/lazNbs6ChUNfcOHTgQuNSoZfHBVHxDPORMviKi0Ku6R5jDnm0IYoNxeSM+U8sjFO
ao0mGd75hK1nzlahnFO9gg99ZUG4GCfd85zAuw0uUvu4QTfvId4wwDFEThfX5fbhlHbi7X2/E1AN
X/4eKVcDtH6NVzV72j0iHli4dvRgZiGz6f3/gUPj9quRYBrrX/Kx+FvgCDseZLewJdLoPtrlkVWK
kZ6CSGd6wnxTva0Vx3aDspvugMkjXt23ndCjozKRq9OLYLb+Y7Bwfnq8Sxm7mtZ4gLYelGBm5NcZ
/m8gPs8oFnpQtO9uE0A6hzeABO6sFe3MLi0BNLpGeY5oagpxVeof/e0oL1m/qGtiAnKLtLoU4pB6
k9nzzi8eQgHZxcJYJUILoJbifVXMg4BlqBl35cRd9uBEbNwoPTPnTCZen1vMBXcCpAwer+2xbSZb
R5cby+SK8WRk2jkcGYjk65LV/tCPr+RrmLeam2P8ReBJM60wq7/LtxgHf7OR7h43SG8Qo+mm6tvv
Nq74aYkYgwM8f20OQLevaqvLbwdtigeBMK74aqQw7mRF38bIlVtYqafEyiOjy7M3cjmB1WqT02pB
rYag82XYmsQDn5kCTERCPo6TmvLeUzrr0x6UKeZzGKk81FU+EewwLITm6HXXQgQIxNrV2fpXQ9K2
wfLwJISPqInTLKrhv0igWuyVXC2NGPPLDdfA2EUqxRNPjIV92gE+p4psFw1ujiQWS1vMYUBXf7ny
j/q9ru02pzYHp63W1HYSGo3yukLWq9HmPybLL4uB7OKV9nJ2Cv/JhX2zwC29A/dCWNexduRmuW6y
ky24VFWuaX76LNEi/3GTHeEXg/435lzGms5zkvarzJOpkMB/VKwZl86eslNIYwKCSM6dMtRyDRcV
HD161XVi6t/ONgXoo7RV0RUyJqVyAEhhAmHamvsu8roDtrI717sDA1SCvo+k0+lZZe2XymARv9hk
ssEHjsvz2EcDbc/emtJlhsq8nf9HNkMmRtzZG94xoHsfKsWnI3T7bBTgEbNBsmfi7MC/pTnQubiT
9lPMq6FWRsJ3CnmEeUIvlPX5mZY+SfqCm3h1B07manQdqblbMFfD/e1FlzogybsVP+RimaN5eaNR
P3yYaqq//IYXNVvqYezuzlsqUg3KiHFX1vETZbnHbRxXEPdCRJJ8Ms4JVNofkOqUAMdfqRL8syQo
ojuIicbJdKMSYJbI16MKaDFAKYJx1/AHAWsEkgVmgcF4/IvRUlXgSL2fppOTo2+TR+00i/2MzdO9
dln+e0wxY802rTgvAa+cD471H8nxf6RlBJfvcq1yJzwd7mQJaAob9uQVfhwifEDIXA3XGvWJ34Rz
F2WyK2kId1duo9GB0BIPzkj800juAqP44BxzF7j6xdEGh40zLdr4uVomUBbpi5+SF8u9R5mxWFL0
5NYQMH/2tUT2Hr6J1kqbPW5EaRQe4ufsOqdVth/au23ZSFvVXJh940fxyavmjhelNRMLd531SmWf
ZGQhCIkvS3p2kTU2f7CdYT7VKY85QRbxTh1NapSfkEJ0S7V9FB0f1b3UxridOyEJBDD3A6QQ9UIX
ZtgkY78kQzB8mBqQ873/rE4pex5RJLS/pIOzEH8H8t5WGfZFzvLrQWADvervXm6Qw9UUB0S60szO
1J2awnFmjI5F4Vr0DenaoIXuqX8CBbrvWuEtJwwvNMjhuQwuaxpH0D2e2LRmGxSxnY+yGUsiCxZq
Tl69YoVlqceU7xJSDjD12zdpMspxsx4ndvMjkvckwVkF2gf3JqtdDwkAIG71Qc/YlXrIUej/jxy4
cpSRw6XOh1b43kvv/I+QWOLlxt65B4MDjTquYSX9BrCyZ+njAjjxE4hQ48QjKkrY+HtO3O2i3PgY
4MGhsUrAb1Ef8kijAGaQhyyRKwgBEfXdEL0J8tmEAz2Bt5h4n4FNhLMyE8RC7A4cJIyDkhXX888m
vIVuXEzQ5xPjTb9TQA0iQ8oM3v8znWcbZHGixwmuTjvut7UUJsdKwoGdzemZtl01fH5vCidmtZRF
yhL2s9xFYYVWj91djbABRfRqRPIiRQp9MUyDjtetFBED1AtWZxsscEWRO3+OnjtJhZ1Jlo7vldPC
qbj9TRVIJHxx67cfgQvBYWkigzrmlb+pxucd/dpZLI/asTRf1aZ0U+qGo9Q8fUPr28M1kv/63S6Y
IaLPmGlyWOkrDqqYsMTJJKoNYYM8z60rf4n+x+nheukToN2rk5r8bOVf3wfQrZI5WWwZPTWOOney
vPmJfbhk/xEnnRnl9bPyjOyExMHGnegIbm+hqpNae2SRSVCz5++J2UZVD757bOafb9+KIq28MqrQ
pYTnrJNklCPZbL1WIRJ23ry6Nzm1rcngXflWgon4K2rnE87VfdQb6mDJZB6zdH8gcwzsFmORqa+6
64xsTwjNCLMBWYp56TwB2h6+yTohBcNpgHs2CLsoVCj0l0NlLKSbTWADwW+q8+0Wr9NZcP06f9Dw
IOm41F/8LiDaIVi37nt+wATrwGsfFa0MeHZoE4rh128QkoHJfXr7cQWZTnvgB1NHQ4A4IAmXhgJ4
xqqnoG/wWQCTMg3s6VKyQzz9/WtbgTKK7RLIhtdf7zvqsp0k9aOTAlfwYOAmEZm/v8OykKxLi+CD
KyvvhOLnKCS0pCZ6tQNUZdnWbJYcE6RHI7+S5ywDJ0qFlv54+7hrJg4NCz7NytNajn9j6T0Alp2z
vrLwLQo4R+bCbTkXQ6xOdp4ULbH5j/kQQ5y45IYj2UUARWYhR3bkT4F5nmbdfVPybgNW0kruHY24
AMOwcCmsSRnmJB5ZxYxVrVgyaLnAHNvLEunFhkwdhiOhSPUqJFcS4Dt7l6o3kQHkSs4CzBvpAODs
DbXTjWonyPawcjk2ZmRrTGLKZ1ZeFJbjSljGvnWDeZcKT6beoas4Fm0bQCJ0jQYEKgRCIm4xiHYf
jgLqEMMVqcZc2KTnZ46kkloxY83uOEqgOGhfb5w+z+A+PvJg9zVC58/I+7zCNnX0TqWo9QAeZN2F
gl5QcJVI/QmHxDP57VJnBRS9BYw7nnI8SBLc5XCLbprEUOP6fUd8BEC94yRuvJI2nQPQWstNnTwr
e2YGmSY9OBtqI8B70xJXLhajiSWmJ1MVCk+UnH/BKYDNrz6R+A3+xNNUDGwLIb3i0WLO1TEhG3tj
Nysfgp/PdoyXNPA6o7mqx8fsjpnCWsenp/n6aQ4zXIY0a90zUWfzxGkRZ48BrZTr1QSq/8SCQDsu
sd8SAKowHqAIw9mVQyafyZWnoNmT7ufWszoMGDT0tRQMPH+8vzEkD7ZDosR22231acGozoASbspl
L4dPf9xTBcGqzT1S8bBWvcmY18BjGZmJhyYEJpABLaiMJiASEgbcvQHKFffb3r5f+dEiiI9pUxAT
jeGbEm+nuw5Y9bYRj1Icp3vrogFk9ou22a1VZm2+79mnRgDm3T9HCpFNLe1maLklJxqH/A1SBReD
PrNEPMiXATnVZ3uJpf6aH/lY+/9Iz/99AhjBD9h2DgPgUkXqFK/xcZPRrFFpxaFu761CRsk5IwOU
jPFp10HYzqYMLBWzdaQ2RB+PZfISSlD50kPU6qnh8VdRUgcZbSdnresNFDwHyVGOmcIJVwkpdR4H
dOvQbAJw2X29DlJi6eSj1hDM1uHzOuWcATeoYqvzgIkEu8JfUGheUmf0kHLwGOTgm2QpJOjeHHJg
YTM11tg0AzJRqfWdKkbowwjgyQjIB88Vush93B8wHNVhnOtETZlKQHghcqpwp1cbf44VaPu2C9Eh
vc5mC+nriTYgaXKzTb+CmhYi6cmoAmB1EGrvO95XXrL43POUenzOa17Rjwtt/PY4JxBBhTRmoECU
ESyfyYABa2WejChF9a7tFf1VsluyY1akLInmzCBCyLkij/qUhG3HtbhvNnfNjDFgVWlRqA14Z9Kr
tqoRsNXfYlpreNeQHN4lmTXyDEMxObBhbPggD9sWYTNZZotX6oNTV4uS1eDh9FFACAF9r1+9oaxd
rb05k1j9VLLLAoegpWGcuVgqT6CSCivsaqJIQyxCqA8MPKnNLUpsGVFW+LnLZTIajqJe05n3EGPi
DMJotmpLxRvgE9LbSHrbCaXDZf1pEyj+JP+NmEn/61hK/+7veWBECnrf6nzjTeK9n3dPmgDbg02N
7sLsGo6iK8jKnXjIIfL1hR/OYz0Fwt2ZmW8qDuguA+NmGgr4ThwHeKeoHoBp99HapnUxlFTjHs1W
w+orGz6iUzAcGQU/6NT4sR+VH0yRPAAffeBX2ITBHF7or/MMohRg7jjF0Bw4okQzk/SbJD4xqBjU
LgwG/jt6wpaoHTxD+gvAD3ZlJTqqz9DKVhHC2EyEixKM+WKFQ3mFW8sZB2WYJ/YBf3a34NkkO8k1
BSoq51tJBhDhS1HynT5lbHX7KksAgzuVUolT+uLJYi41AhAqv/WJx3/kUYFnBPPOz8c8HSfvK10d
tpaWfu7GgIe3TUP/RHIL3Y+CKvzmO9yJCD800GlD35pKVOTcQImkmiN5iMGjVzlAFRBXE8HqDdxM
KlU1mlMY8R6PREy2x93FkUx2wBZbU2i3YRTeyrEIADGGZAfsJ+KTC0J+jUr/VlaECVbtTARoWT9j
bBv8+A+hxfRnK1l26NEB1OyGvQ4xTPrR+QrtWiPwq0lpzfC6kBDfG83IBHD/MZ/NfT1M625nQR5O
0LliKqHB4AJXixgFPfpmyeE0FDCllm752P2zGsKe1uIXBXa2mcYQ0eonedeLfA9HoVbWqpSno2b2
yLqm/L+mI7kVmBoIG7X6DKjDSBkWUU/wt7k8OCW/bdphh7Jx5XIMzUMmk0DJbfNwW/Jiq4pAMcHB
3GQRjl3B1Tn2LUfH1KH8gjoqqH3R/QXxlqj+fgwI7mcfDAWTJS32cKmcSsqDuRMm7F3OIZF2PM9u
/enjPjeJSmh+Z1DTevjRAQx7BIqYmRveuGsCF6q0EKX+wCiDkXXMCyvmUHRrrKMYgW007JDX63Kx
Bm565EH7h52vjvyiSBQVZwn8GUWPKyOmV8W6veBZAF0IHmyGjX95c+9MrMNY86RDg/dtzjyVw5Vg
dfG1xP7CRp++k2vLLTQFq8AORwwJz5dyUkr3occvwTzbwEhUR8n7Bm1QY1Ox4wcPY5DcvyiePYon
shM/dfTuK0MtZtZvhPKuKdn6bwJciw6ymAryuSO0Ebc9IvByMMuRs/XmKgifWffSzms1ruGyYvT5
SWxYZ7XWt4pJYkcT6MUTwfxG6r+q+bV6LOSxeazpZeUKuhXDR6YRU0WYA4nFj/8j6lIUAZ4YEjBS
tHinwEx0nZDN5TNM9ePW7ZmnGX92SRB5yoEDPk4/SCLwuXK3acJ415VLo7FoPqpjWz12W9bdJNBb
mUQiCnHu1RpebinMkTV3CXlddEHx/bh/v+L1EE3805+vl3Hz2HzIt72zZZJ3Z3KnkpBhU+BzAlFv
4/E1oDple78nchOMBqojDu6/Mfula55OZjOeMOGVGQgBgZsWCpQxb7Y89UmqWT56/EKOOtoYTEFe
xUpN1ttw7d/EB8nsTBN5asN5XDgft4Ky7mFcmLJcU4zoV4+LyTRO+mI3VBzd1bQlIgYzl289zQ3s
C60uXyroLwCRsy8TJA1Gq7fcjzMTDawkieai8WWK3rlezJyr+C8We2raHDYZXy5KNDNcCjdMwmXp
8jbNCdML7vFdxUd2JfYQJ2UOYeZDOEMZCQrfB9b7+qA9AgCWuq9PTx0nw4eOLR5EV8X0/5wG6Pbs
Pt6zszrEWsjXxepKtJEp6WE6u98WY0h1ArW+dG2lMBHO7dlg0smhFRhZWQemzQttJuOaGp/lS7aR
RHOAmzZJiAsST4MB5mK0eIfTyZUC8ppaXxwzg97o3Y+yMwS1OEASjK0h7TJMqmhtZF/p/8d297Jk
XOK/PvvWd3gzn9zBKP89f8c0D3lBkqrBC58HGKOLbPB+bQlTkXNnXM3cuobCogiR63X4LrsHwELT
y9AxgqOtGZRGAUlCeAvrTZpI5PZ4CwdrU4853/ut8g+w3/vcqcWno+oGm2DIAC2Jl2CCwY7chrF9
auqLu88dbc9THRzqe8m7hp8ywOw4XdZ4Dvg5YxZ69jJCL7JUzLFzKgNQzcZaj35OGeq9bX5mJYG7
QR1G/IowooQ8mg1Fdk/BsrQOGKdG2zxxBI8tbhwl0ETyjfECxIcMVkkzMoGZUmYUNzMJooixAcph
Zspx5d6O84is5kYU/L3GdN4DMJaDtXYn7CEHgAAoWttZGwI6X9If+FANicj/zsjtZhQgt5tYLhu8
1igQopjJXdf1ybEEAwN8gTEtGNH7S02KvdaZ21fwAkEGlELb/o0DQU3/TEgWHM0bMGShHdPRuVLD
IOZjAPkgeGli0MSM/68wdz5v1JqoQDGuDd252Zl+gEF29tNTCA9yslhXMYU5NhdHeH5QD7kU9dcK
hbMAIaEiIf7OWaVKZPJuHTvXTvfn0n7ezLdQZwFVCGDDTJfhT57dS4Qufq9UMKtLymaEI9l3hMSv
ryTSTF7/UHB0HNwougWQ1Vj3f3B/F2v1Pj/XNxxuON6CnuH9/bnkpdJM4Mh14RjPGiDyUrL/IM78
AJ/cxuSYSk/UY26zdjAmnJMjlE2w1TMtM7SIi9PPzEj57aRzOgU7G/s/t774UAmAklG2cbxxYken
VCAE/W5xIqWlEi6/t2aJaLh66WNK9i1Vva6IGDQr9aRCpvS5ZnlaxsQIfOyb6dXHVCqZkZUYdnxD
+xvwnyU/TwXW58ukgezmvjCfjRbE9jsENRPlCNZGhoZ8wOz74J60Xls9QG/zguwAL0VPT63p/4Hi
BVAwCQiYmyCsWnRQeMMVPhPUj1RbhdK88biLSbT+ZfuhTLbFluiXP8CCum3/kurWd1030TCTB5go
5DPgMn1SedKvsiZb6se8miSBB8cTUzkzQ9vvteoKUmObWtGV87udrprGXrdyG5bOKAl04ZVrKbiB
7Zwg3MN1E69XdQ999IQL878X90EjdqvA531UK6flPK8yvE9m1yN2ZupBgxwDJ4UFOLSOapVk4hei
BAjpeP5VmhFje1+PyZzGkmPgVeB0tGUjPa60z9e7pO7I1/bI4Fi/rwY0HOo8PL6afnCGfvt0QAcx
HMGDg+QzYwgwH09HyX8aeOUTabBBlgHDf4z94B5P004EfH4xhvj+/uyU5SKdPgDNNUivuT3bPmwv
VqImXq9wdrVID4DWX40uUlAK8m6WM5zqgU0acIqLMimns8gPiHGptUwBhTRYapFoBfRrZ+SqKqer
N7uswptXD/M2iQHuoboD+J7SvIRpRrdW5nxSZJ8SQsgNjQ5kjqeYPmnoQ6q/qJzz2LVThxuPwwJV
4dGUMs9TyEEeFy1y7rWUgQMQiItmLjvBj37CZzFFbWj6fRsDXzvuK6rV+O0HggZZkMaiIx1seFMQ
u0Kvd2YX69O41YWGZkwFAllDkzO1wGxaSCWehjf/ruA1xFyUqfExl/vRyYTAM6848sdV4svNfi/L
G0qZEaHF/aF2HFPe20CxWYvA9CVlKFnd1wE1E3WmeFt6G/5TQvog6Egik+oAQxVg1X1Vfk6eE+Ot
zVGdqs+TvRh04IlG1JYG9aKAVGxMY0ZeSGcv638qsbyriCaql1i3BPCj2qwzWvBnMagaLLdyVem8
EUWVtRc9wJ2+g9P/cmyV+qiXb55jeBifoUVVxbHKl7Cl/vKJ51bltlVpBy8iXr18Zvhu74ivvfc7
Gu4pjnrbD+8SKet8yJVrF1BDhEqC72I4icbZJQuA1hI5arE9Usoft/sD7QRyjEue0nzlteSKj9H8
NtBWtT7pfQWPNKyf1+p2t7Reji/8AUSm/uqLUPIs5JT/I9ixdirOqQsi93fCEpP77X/PG8XoXyGw
iZcWKaG3T8MyvibUXX9dBeUHS4C3twIl5+ogiUTImV1WYVvXhIXEdrEI+iYqn8FCo01ydR3ayc0i
BReH12V2jGBlXhz6EkgVVZ//UCxxf2rHD8wrY57KEwx1zxHymwT2LLaeHmFQrUaIXx161NaWKMDH
Q9cF1sRLwTgPMasvFJwwL+r9GqObJZEBfVspoipG0iSQSy+bpXIpLTHWbdhFxNTE6JPADsgMjJzA
KU+syK58NUqaxTKdYlCAoqtivMBdCEyfaZFkaNRWay/JrE6MTUtw1fWLe/t/Aw2J9xGJjTdfNes3
XwfkW6DNsszeKlM9USsXQVYqalHRjB9GMt0e/uPpCOmNM8shfYpCxeG7QH0qJUG+Z6oMIWdwx+1Y
x5zMrsUcfXvakNXFERPSd6JeAPw35xyl09auNe9+H+TKwqyYxiTlawEhyrUqAWycafEY+oEFRxBq
rm+8f7GE/4hPFVy/no3QFZbQhtzPtJ8ZQvm2d5w/N60g99yUwcxEh/A67ZH9sfFo3sSb0mv1JIVf
Gf5AoZFfeEDVCY/nHsUrIZornCm45R8rt+GBmO2KU1lAQOFZ4lzWkc9Km4ZyRuUNZbcZscZh7M9a
NlyGzawHunqZKiKkVeMMhmsKpsa5bhMwgOWtWcTj4P0LsQl1TNTLogbs82B+p2xQS4zBwAlmnCCT
nkOpIaYj9BL5J8LxFxquOl7ZlSMt2UZSGFdFwMjf7k55atUsEccDYkqH0ybTbOpzcCMfZx4Lkn8B
ctL8YJt4xfVwYEeykxwN2yA1gnIiPsjWG7tPGe45J7/diqnkQZpwFWV0U2HTdka5CjLx4Tx9OeqG
SoSxKu41Z5JcTUmwdZ01e0m8eLgGtu3Ng9yjRIueRGsYASf18DRuWFDO/lkgAvw+W2xrixXhm2vX
BNahA3RNnVXtqDTuTU5qFB08uMoabdArbNJ8aA4+TWsxqOmRmnjp1E3fU808lXi5Q4Qxk1mHrL3+
sU/dEyVhx9sOPG/59uCEJbPOWdMjPUomkhit6e3qnFeeeVz/kWW/6pBFGXeiaXKAZLl7prK5ZL6T
5Wy28WnANyrpQXAXVkoFCWzYfDKluxMlbW80/WeoUiVATbPtyACSdzDoPzVEa0NFFGxJ8x3NsR+i
JLmA1Qknai69+f5DDq0vgr8QJ9DzD8xBfrIoHeuS+xjJadpcOIEDJyKMQRr5G/SYlmc8JggRDfiX
ulQG8BxUFjxAdYO93ABBYyJj3/CeBsVg+Pi6lbJinfyJ1O8ABeTmo3yFDbaMMj+kNBQ7iIyOnIgB
J1fG9BTmWQlj237L9+HOV7znvMDW918Dsir9y6S0elocW1HQ1a04gBbraMZ2yQVXkewDLvgMZo0g
POnq9caOnrh0I5jzvYxO/66KAqlCEMBFh4qw2DzfGNUguhM3rDRdLnA70DrmSRHhMjIwO95ilSxR
FhcgkwpWf5NV6tPud6DIhPODYbSlJn0kv2eqR8NnA+pRHjoa2pFL+18lV/GVYPC6xPSlYB8ESZo6
TipSITgzknsIQ9E4VBvzoeiIzcgZcJaJ9x71HkMgsYiW8S21FzU8BF0+GjEnfS7KGPivfIWbetla
WDlpWtSCCpoHMwSixLETr5Me+yKYyRq1LQZ10Te9+cC/EhwKa4g7i8huQ+KGHIyswjaog+9M0Q3S
Xx31z2VrM6MZ3dKzWSiSLkjBtewdGa7bcFnlJSwzUDhx5fBwulzOd8IQSonOLWOzMQEDA6dN43+9
zq2Q5WEzEQiy20YttPcfsN+0CqBw41AMBVyaOgi1uwIt6I+nFFrrOSePztmrq1yqZSIcqsWbY4j8
dYxOHTnMdy8jvOgOo8nYKD/r3hY6woAB4kp2hOK7RJmdZr7Tus1i8BJElNfz9Nev9tm+vCjZazwH
R5XeecFdxajSogddLvgKlqEbhw+E3smBbo7lzNCy/kHFIPNt+1g7CI60xyAp+ohmudDjqd83CfU0
78hQp7FDxZDjMrBAJvVnyxoapDg/e2yRMWA99BgRt2HLonJHFYJutx3LNw8ulLdFp47A9s9UZwIX
0xwZx8d9GzUCBOhDo/foTg6sS/hNrP80ebOBNOzINwZiDlUD4ayXSQek8RRVmEjoKqGsXBLEYpzm
PkSwy3OIPYLxXsPVwI350v+mTpI3mU80F/cuY9k/PZbh1sHmPz2UjC2DMOLxHm3M49q3+XHrOnUi
b8biKHPILAiBXZJdTGRniqD7LH8A96Yfn00guw3RtW5bt8MLHtZ+WowNd5UF018jPpGIOxBhPxY6
0yRasi52JZCUtTLo1/xHFbcgOjUAG+r2hrzrHJA3Y16nI5rJNnuGAqSzEYEzJ2Lw7TBHLzGHuytD
9Gn6NiqwffGSKZs8xvVbRcQkcS3PrdhrJDzVHrR/BfnK+jKedMQqLG3GqZ2Os65SNqSeuniWjnly
TfFH/4BAGeiLcBA/qD/O6gD12y9jspTKb5A5EKpGZNj8uI7iiU39aa3PEATNz269FGdH6LOz0YYQ
K9glfx3jXTt1I79ezPX2IaP5GUFLLeDoVn+vFmy6jAKzwE4GXV9VeXrL6kWXHkIKMkRdRsSvZLkN
xmDN82HOk/Wf45/nzoKQHx3W+ICfTd+Sgt8apRK/BfcZfR7VOd8Etq+vHGxw8idPX1dz0H903UDZ
QcQUmcWNa8vwi+AdOWCyCBPromXnqJPC4JWHSGoaCg7n8/8NWLhu7Y+hqJXByljlw0PEKzO73eKV
gpGQjJfFW4QK8iOau87RHhwuPBnFOIXJeD4xX6goE7rnzZ1YoB4FmT+vTLIUJAdXWWZXPiCrLnXK
Gq4T3JvtnicO13KjCK+eprbfmJKonA6LHaWugycTgAK5NKh4DKsbKARQTGRBAqQ6clQLOQaOM0cE
M7+z1lzTqLMFZFaB/Wvi9DLSTYUzVGtBFe47FqN+5wRD9UmKKmFhP9lhVgxz9xDFI102CzTwjZ2k
DHDV/bjV4BxL0FQ2mn3R46rzSbkx5yy5oreG0NzGvKFMJ7X5Nd0sQane/vkJFgryArIGP3My6gLd
+HmDU0x1rSN9+OvuMTgkP+2n4rts68+z0QfoDuqCEVYhIO00OBU37vqdPHLRx0ZinVjxWDbBxHKo
IXVNpinQuJ8Tab2fMdNBpzQWlgXMpMjXxoMStV4zPtIoQFSrbsuO0VlFnAUbzj0CJGZef3EMHuh5
FVZVwRyNF9V4bGIhQvgnX0FzYBfFenGN5l4GFj8d/SNWbyiwaCLop/BJe4jvuMBxITC57HgHzIrG
DvYyFHnsH7MDJ3oOpBfi2UBoRJr7ZM7+k9QeeWuNy96J18zUfKdmrGyEMi0+enVeVnkvhlo/6Lh/
+7Y6wozwlNV9i5AVqC0zjDntniM2pxvYt3btLBkkdgL+8ESP7wyzc3JdNaw0mHH79u7+nnSFr0tp
yeQ5g5MKzqJL1wvR5GuCJ/ebUWVAQ5snHJkyyJnxdprMqeJP5hhOE0xawHVkEt8fG7gxq9fNo1BM
LAU0p9ODYhhJzBmVfEZuYbgp7bQBX/LOh/igmK0dbhAoeE1XdJFlG0rDlAAb3x/8LW1McbHGfxfr
hLzsTRoI4l8y13EuWsWjE36StSKm/4NVIY73e7pVaUkERteGBEC5Yo8hL/Jqqgcy7BFnViHJ8Ez4
cV03frSGmBDzEDtYWSkZMpzB5Eu4cRdOqRorFwYWBBtXx93h81lPFCtidynlGfo9GAkXaYq2jGAY
HGQ5ET9mPGh4fiB8cx8OzdjtDkz/w5Gp6wpWKyCp1C6M2p9gC85ElFwNMPo+RdbPEWDLwckQ4Ywp
IAKF4w1dToYER+e1cF6BpkhWFhj55cVWe699xkkS+v6nDAOvcmmVa9FzLPTTjaSOpBUVhmKhr9i/
GLUzQFUSr8oKf7YUZgN/1V2bdWgGXRBrMh9F+35l6jYgVI61lumU452rhBUrROInpql3XsCgByDP
P7yopSJsZ53zr9Ivce2+anGYeo+PVXBg5gGAL4oIAuWEywHFd8Ww8mM3aYgne3M9y4RLVCJq0vcl
Sgv+yuCwMwtfOnu+8JH1s24/+zW9UQRDqpXRKQaKA7BmsXXm5h7uVqTzZTAJrFCh6OBrRgQx/ekH
5wePAk2oH7NkNf8gXwmaZwRUwEghZqD1wIOwGQFzNeHNLvvULmqclSKnMVl7GB+fjOF5VoxX0+Un
+dxLtVGeK4BgnPuQH8hCNncn2ctj8dwjeQDdrBgs8rNmxPVGq05Ekq1WoutyOgVPff5K5K6qxOl3
fpbQVUWhXwpGc8XmgaOOwi14fmeNHuR51h2a4OchSDr+4A9wkcLatO3uCiN+cTMJCS6KoDE5OpRr
FKxffBgNXl9AVm5Qy7ykqI/pIhwTuVRuz2Govgjg37agKdge4Psqorzt4nRHM7BfwrtPWcFkBgHs
ZUuKjAFqvU4vkq/X19HtmhrgSHjgQJeM7HK63iyZbJaR9ylByeTnvMty8BXpmWG7sxutBw7X9Vki
q9RQ9aO4xqXPWCLmLcVZMBGylXU/AhdxxusNTzBmmv/BdGKQn7V/pB6m9/63p/ODDctCBthZ/12C
hAHd1524ek4TiBNkRd8uwrec/Xu68EbhPS/qgXZnCbVbssDXh1I5k+bswhqLthLWEaWVhVC7J1wh
SUPaIusvsbx5u0Soi8Gy/OcsdYqi3ZNWvzvnp9Gy8BNIP4RTx2Kj83/u7v00E6977vGZYUuDlitf
+ohNa2GbJHD5ybHdthqSWy/K0HQ4gUedxbYYwA4NCT43D6CnCq9XbeUyuD6WFlBDYH0Kx4jJs2uY
gRzPPwV3B2F4fAdcjbqO7mI1lrAwg4vliovlkxHXXRJLALwKL4x/XJDhFjtNum+1pE9MKcrvqesQ
IuJF48wAZvgQU3JweAt3sp8y/NiLDRqj1xLR9iY0gY7MMv8pJH/RTB5zQSa399X49otrNxJcviLt
45zXxQsy35Kz5Ng9V2F2uZm8oeit8/jBvR78WXyFuUw5wWtOBOow3rEFjBSge28JuCBTFrgn6UPn
uDs+Lk/eH+JKBabWTUhaFOwFEQWFM4lXqg7AjxSUuk4Sx0lM947Rmi7g5hNy1MeYKkc4XQBMLaGG
YTvA3oDNq/ASOZbFEmC+eIKnFVFBaGmZ975S2KlGQ33vjikLFFTb0f85bD06WIgIzby6XdEDdtuh
EDep2B/b3FIlAz9KpnTWOZ14EQFq7GdzbbcOupDkt89dN8OxYRwCBLWT2sTPc/UMOxtKVhXvjc6W
6PJxyxgRyF3ofpuUguDpZmqRmqAPrG40LQoSOTSZT0wpyRZ9CW+3B2WsjJgOFNViFy4Wv8YT7jMJ
oZu9qTwZ5P5dGlGnMw+D5ZNSRd0fnrdrSvJwEZSyCpJMX/i6phDQV8icL6o/PObc2cdhfrCBsNcR
H3bU//bJH75qKC/oNgW67XedJN2G6QwBobheK76/jXvpcU+RbZt2BQ2DI1POzjpOBjqp+gL7i0b/
ZD9RdELLr4q8Cx1cUaVJIqGwanQqGoaJ3BPFlOPouNGeBtjUchDUFbyLI7CArQqYjrs5yeVtHM2v
ERB7NiJ7SMXWklykvtX0FsFpm9F+mw9TnVPre7g+yHmnovnXw2BFgLFVmxenoR50H8TxrajlzG51
Ia+BhlvULl0Vj0sLGQi4KQbU/nM8fF+4bSYKN+qEp/UVIYvVdAXHhSS80eLvbQom3kGjNyEOB+7n
1kQ37nSCkaWMOgfIexDp9uOuIPUxZGngURhFYFHRw/mPuC17kdnKMGGfII76HCtf2Cudxpx4jm37
8BP7aYHmepwaW9VQOsNot4dIRcDXWf00+nAj3nSoIUcWK7sBxuH4xlcMQCyWVxomYaVp9I49inDi
eRCOJQAHXBDSaXoJLNdf1X5nPlp61KORJcGbwENQLucuXNkD3Mzdi6Igl/ZOFwgZ3m0WbVdJA6if
AHMkjLlyz4QYIbhivEcKGCcIgH1j4ylLdwq6e7uwKPcM35axViwj+LUtHFXBRdGum8NaS1GQdKV/
kNg2CgVoBqr0rQvzRyokO7NWio4xdl4PjS5X9jx0niJO0tcKmkMx8mwhuL7MZ63Z1OooggxhefDa
mUxGQfdqnQycWeAOTnnNC5nRmjYuNO8a1cwySBWJZupXufCouJBkt24gOq9xDYpYSwIp294boajK
E9wFBEs8GMxUK26cGyBUgD3FXwcO6Ai30L3mV4YYXpcsKNtsseV8Rmy2DZglUAek80C0Zyzwoug/
0+HJTWqg4GtBwXclnXahozPpGyatmk3zYeYnmr5wcLCdQ7rs+IOOKqMXcE67UbZ2ztp2r84A7/mo
5tmHy6py3yr9GBuYWsDDKdu4PJ+wxokhCxeAGqKA+jjHo4FJ0iEulyLTh980xpeyo8JsFsrqsHXW
ZLuV7vY+0U/nspykKUHzb4AzB1wjjYt76ep5MamEBXRB3nJqWVt8BjjU2/1fv87QXgiDi4FaSCFZ
yNVvsyUBr8cMd5AMlkWRuhJl6QFyNZpRGelmzkeQlbkr+c+eKWbFWFPznPYQ7AG3bJz/gFMFIxDZ
RoVdZEGYDCvvIICRYnbU41kRAKpa3zxFs6mpZpiHyndWNIwV8cB/uWDn6p3mfFjLTespO8JOXT2A
XKMFQd6ZCzU5fDGl5a9P+EC8FlFCPbb7RCk2N8JZxfpETiV1SemH0UtophwTZiLfhZjSehe2CxLm
m25lYot7qWpeMtxZ+fgzSKlyp90UZH3wnfUyMvebpwnB+FVU6lnH9whTDyLSa9Deg9O9DbpWPSZe
Ys9OPSMfjERc2sPHMKpzmzGKKBHaFOXFL3C0Vi2KPKj6n17o+zKDk1CGfjF7+NuEf9SCqJVdSZ3M
rOFIMpO2Ys7HM2tDGThrvAPaKw5mMGRN8ml9czM1ECbLAbMbpRFkvnP93osULgfJ9hpKPIydwMCA
59Ysat96fWYxxU2N6HZlFcygN99obGX5sqVCJ1ICceXW2a6lWX8qxd06G1/wfU9PZpAwt/ouB8+C
fyrJ1YoMF+G1nxuMDsACpXzGDTij9E7Myk9w9PXWE4gGx58yr8PoHF3oUomhexK0kyVczcmvd5Kf
WCwBvN746TyRTk482YHU5lM3AR2ry1zM2YStNksT4FV8XMWmZXNkSaAdef1k7Wqoo42FnsGMK2KK
xFtraCqOaDzarkLi/Mw8cscE2w6P7Tzkp59vmFJbL4SYVgBeNk96R0ho0hTMUMwoL0zxut58uqXm
rVidI3exgyHIyQQ9Z8MQ5B72IBlAZh60TUjFI1/d82SJ2x/FQMzyQCCU638hJ82j5ZXOe+DVEvgA
Aq8CWlvYhcq42alExZ8IpV+joSmMthynLyxPzPEjYvjEx+AWaqdDiGfRXbdhqtaj12uyrhbuOX59
PJ+Mo45jBDsYXSFPEyBQ1BazsSu068ZMzkz9SixuuD0hOlIwGB7hKyV2Av39scTIN4VyZ0iuhuu+
ew86fsDGWLPOejPLoyFhjcxOJ+ntxQzUjnY0tgexffmV1/spxG3hW/Adnq7R7+L2fMD1SxdtcvZE
wFzwHsm2INH3BHdgkadDvopkCfTje8QR9IxDsW+JeyUAG9vwcS99uE5cdy3wSBoJ859QxnAM2Y39
3xePapKgtDrpj9IlQYN93Wh8RWOUky+7rqf62KO43b/R+fJ6TowsQ+7ZIwedziqQBIQ1QlYDikmp
KMsonIRdNFuW6oYTDp7OJa112RDBgcsfewkUPdivzIB9oBbyA6Jecf20sgQGSVi3zMRK97oCLHAv
ELOH2W5s9gvboaRgsoM4eBq/FSJkInPGkzpoxzNy5nPfQk97vw7vg/uxddiGa85yhGlTKg7QPgKh
3EunZnFa+9v8TmHvsSuDxIiQtFiDLz4b20g9Zca+mNSpqYLyRWSZpNo6EVV7qnJR+BQBwBCQ4Xkp
8UcNQhKzAWsn7u5+/19XZ4itzzrrySHyodL0zd3xcf2451FERzn6LUCMugkH7NUuOm0TxeT1QxeF
mhiRLcaIBlELd8hCKHhwOQ+X4ayCNpPA8psfpZVi6Ayxuba0D74rW6m1yNhwNJtIQvmb9b38AtZq
PBnZWV+n4YWviBEmZs81pJzeKz4+okO2Mo2x8e02A1dp4RFYOlRUW0wLC3oKE58QvEbxiMsIyEb2
g/bVu1wnoOTWjCZ2T4XOtFclSH6iMv3NkXmteIqP3u0Q2/gytNBL8IuUWr7zwxAAewxCSD5UFKUF
vtU+GC7ySw7XCs9/Os3UhUvctJyrQoG8i6BNLzoxSOhcpv+YCRwP+2XMSFoXj2MnC8jZ0OOwPCK+
RT8fxMQm2OWOjcgYIaujZZxrD3gwY8uhAop0LFAmLJdr3oFMwtK5xDcDfmY6s0GO6iSZnMYHb2iD
KAUWXBuLfvx8bBHZ5aG+DdzlcImyUyxHmbsPU3fTMOPOFi+/EGjw+Xka39hhlBUndheP3JgrvBAe
MPL3WNLZL/1IDIGIOFBljpKeC34B/fdz/dm+3vonZS+D5AhvILlSveOEq9TNBDGWb/elKtpLegd6
P4RUyNnN0Y5x0/gdW4Siiap1MuOkDPciDF7WrCWZOhFtfkMdqyg87+g8YE+uzPLzpS7pBxTqZKp6
d2oB/9zOZHldFVpqwqH5/TVhbw7X7ybOgqUHK/KaKF8UdLgbJ4aUnkT3ZftRg1TBlU9RaXcn13uk
x64GUmVAWJ+znPMyx45uST7RKLUhUkd6MJyFwwGnrzGuLRgfixHBT2/fYwYMSdbGi+49srQjQFFI
kYcT0PxG2CBvM1uI0rGyxxMWJ275jHcPXNLE6ZKy5NBkvSLdhrKtHyQFoSN+g2jfnczIJolipsgm
9c7rLaHPF3O4qHQTAFOLcAhfPmWQD9tniaWTxFLe+yt4rTSeGB+PADnrDaTsWFAR2o4VfgBibieV
HYBAggsoWEDBWBMF8pdT5Vy1HKIEpREeFnW8qS/+pt/3V0mC7zCa6uS2T+1yOQdKN14GP7vn80uM
u8DlcQNhOSFyvcch6xtoY+00QtFJFshybE/o1iFiC/r9w3TpaH24QNsCLFr/c8aGeSFSCF17nfea
c1Jl/TUd7fAEjLY55nr0TurQMrwrBaf3FGc+dfdE7IVdX80mUyEgcGKmsupHUPyelYvQ/EGyAjic
jGV8zZ0odUvwInu38yFmPnWls84B4iBjCZB8eZUU7jF9nB4AL7D6Uz3guj6Lqhfih4gNmn2lxJuS
2BTebG1hMGWQ1OQhbFfrRaxNhX765vlVwGqTvU+JlZWICDQI3joaRGWzOqe6aF3pvWP7GBT45b0Y
iZYISmqomsBbWMsveZ06zWEkZEGljmyqq7Av5sxhxSHuIzDI8csERJBdzb89y4EkFNWnIXfDQHNc
x9dgja5WN5yOcl2LjVM5N6ZWtASqNR11gSm56+p0lNlyixaZ5PUxNqOZXJtpZnyxq1J7TJX/8T6L
8lxvi9+qgeX2KF2E1jICbdyfg6hNGtUATf8vYhrPWAzTSIwGpUjCnOJdhkl5f+X0vAw5xKLsISlG
7QXNMJa6ztaWXghphY++OIw0SJKgtysHwdNHzywhYDW8mPUX04/SGU7YpVRhiJKAlvV7wy04p7ci
2AQ1cquTHtbnqRbfQF1d47JblCdkNGcYEfCLllK+a1DAmNO2ftQtbG8HX+7bSfGtimDFepakEkGz
OuCaereAUFzLcVobQ0T/KT43r4dA46DoDO9Ff5P5ISrszwQ/Y6EegNPMFRzQx6GeRRJQdsLso8bT
M8grHSgReoRHtkQ7v0Ix+odryBRmoqlEDQzWIYWNfwhj4MVXiCqBG24oUiYziYcsxtVghlzSyUxq
MJmLrEHc7dLIlSCTTiIw1MY14nUTAB/hz6Yqlg4zhALc5GQMj0MiVFpRStnm+O4b6oQWiysw7QX5
EE2ikJFYC/OVimqvLsR+rwScmeJFLOlj9f2pxUmfoimKn4Q3G3viY8Ek9XaeBha4UjPC0X/Kor/Y
+zHPnOko9zLAFbtWm/8ikkzWqE1MXI3z87ACz8H1pFryAHYS3ymXk+qHkImPdiWhTkf9tfFFY9T0
S4jRMlDOE2+2fuNOutnmCnBGIhzknHMQtwuKEifwJFNRGG58YRJAzEaU32x+IiCISDotK+dCF68c
nqn9rdO6L3eKLFmlcYqp6YJKTBCOI3RosOX4QIewZn8oSJXzRd9r2be7WownH/5vznxTrNH5QL4Q
kiVOPSQ1tJ1u1SaKgYsnzl891ulVFrqVrPBSY7Opx40gysE4ZhrUwRYljjf+QITgtWyP4Fewjih1
btaEoJ9Kk/q3E5fhgSg4h8/6/uVUWWoVIPDhYMgEeCP75akXzOKbVLsoPn4R33YohF1zVYsOmX3P
OuGrc3qDJkvbvfVLFE6rPoGyM4XWiKXuJn1UbPwS4UmvucpUAwcfYc7kW8CTSqZjkz+uNdItj/al
3MBB1Rl96t/R4LCpNY3tZPrUlszBOfYA3WXfXolOHiCgmxBZWao52z04MddYAHo0qT+v2nnsaEz8
B1lWnqgpc+Hf9VhxHaqSFON4n0H0sO3P13V+thFGZQdnKF4K1OXCrJgmWFBmwkqqqS1egRtJnyAa
hA1A4D9O0byGdq203GHm7GywQxw9NnVKprnt1XPLqB8zj8X62LL4zXFaV5szUBHWDdVgcR09oGB4
eYl+CGDN6JlzjipRl8wSfEVV96B9yW6gFs3k7oUVtrpzmfBx2MGiXCutmto4sRMGQGjT1q6j34KY
Ouik71wx2mFDY9ee590LpQrTn7/NbXK/aS96ad0xqs/Grh3mhcALImCLTC711WgEkz1yfwyrA4L1
/vo93aAxpsiW50uCF5q7nhaEw6Uh7E8Glo2wc64HbE3dy+otyER5iYOlrGLCBZyNLWXl8LU9H7Vu
JXchycZiq8M4LLLHm/LJJu2Ax5o343xq2hIzKjJWt4ZlsQwvYom1eCYw/txn3U0Z8/eJ1Y7Mn6sY
0QGBS7fQfoFhnAWU50/Z8rL/wF203zzTgCAJMkM1P//ts5G0/Stm13UDiMif6SoOL8Q70xbATaDh
Iz4MNpL95Vp/rMQqrepFIFvEjsA3A+j3jg6fNNJC+RZ6WqzNX/dm0zwINGd1tHNqK8NZLXeIsYgL
xHr/qr3UvqyeqWkIwJMNJxQ4OHvMfFjB66xGo5ikCRwZq+k9hUwybjZJ7c4LjGu0uK4Tj/TseKUq
94YRg6R/zYLd2gfXK6yjlcMN2uK0VCWE7Fegqjxpk3q/28U94kEAYZolq1ilGeMnNoHegTnhAFSL
cBCJqQ8zmxhwqh33pFsebRcRbp9X/yRSmx1aSqdmSB9LYmDt0R1E3IWXlcQGTAcHXnsHyxzelAbO
Kh/T6dmHbK32DHCp2MJf1GjAhfpoeqi/HmPuJ8dEDbZWhxEBWbF+pzqTKkbgfiHsQJB7kAREXabm
MBTdjIleGCd1WuEFL1W49KqIhuGTqxSy0VvPCjLGaD5qufOGgqsvwLFxuYplYW+rPAfdMKjYDF6j
1pUURF5AzNzJPFLjC/1byxg0/yvc143BHGic53Q7mGptSqEqXtqJolz8biYmTYgapj9UyMh3bqr2
Cqz1UEmybwvB/a1gUAYn6NUI24q2Cdwx+S0Y6axsczs2zbcc+yNH//cToyht6vE7rxkO8cyGJq8X
9a4SqhIdRjwPEKlJsleigc1yDJMUXEhZcos16zDEtaUna4ritTAU1EsURZSpST9Sk6B3bueJlYkq
DZurealTb3jOHWZrplIcNvSrLmoCRA0dQpVfqOORI1kbXObpd38zSl5aSnWwV07CYIfebh8ai0wF
GIQM3jlBzXCxjxJ0Q6OR0IfsR1ZemHvMe7TCKlb3FhYlqRuvv2x4mhSAnfLH8O4vSxpCp82+GkuX
LnW+d3VO9L3EPO7xQmvZikMT/T0Ipz/e4T6Xy/PmYigv5h4tHklS7MP7S1jeLpAxIPE/meLTUmxv
LQBIRLlmivL+W6Vc0SncrPq6FvIB/nKANaMTecHU5H5bG9ETD9ogi1G4/9XxW6dC6+gVIpXtvP0t
phegzNSXWCR4rvdDdOMyxd8uMJ3xP8k1Ccg42/Cvv+UJ6PNYVASPrscHu1EbXbaEc1V2A9GqyRZ3
W706N9S+WlOV4OG6zr5j0Odr8M1TJLfthBnK1VkwB+RCfP2THviDY+z4AyWco/3f5pqCO5JR/XHz
WnCTPFB81Rmc9KGoUDllUGFkG7LzNRTA4RDxfBUq8ICZqBaLfNpt1GU1W+fP3vWPbZ/Fklsx4TGV
Rzm25pzO3b09De2b9OT206d5X0Iuun573ZXb49zTNcdQxYCUFVkp6TwI8nrHMZmtNRrZ5XhB8cB7
CMOWsYfZ76eTzxL3Ei3qYdEZJuI5kzpoPnor0ZU/7O1vrdyE3rDYBHZyEJ7sjbvs07NSg2wLRMIb
MR1xTByPm/sVcE7ZYUGkVUWZ1rYnYu2yC32lC3xyEM7V9z6HCZAx5f1qBNVIOgHSUB+SfaYeAShI
y4ph+s8EzUgdsy1+mNXnzc+Q7JMhn4E+p3QlFOGGeY5QCAzYppmR064n0mnbn/cvaajvQOWdbQkX
MBxYrRB1tvJNivQizj5kGDj4M/hoRYlnWMSYXQ8yMt1bK4vQ/VTOYjCncOVlIEj1i2/6OBnNj40o
M5+Hg+Ecbmm8KNNHYpXlQDgBsVhiAFi57rpiGVzYL5zr5985Oou6j4yjVPbF5pf3ZsNxSx1//DdM
+1VB/zFcUSyymTYDV/r2v2fi4vDOH70Tz6WK2VfJGPi9WmN1zV1/y2R4GGD6ATp8BULXHzdVn7RZ
7KX8s3jvB345AJyEJaYFxwCVVSYjGJ7PtvUvEjktZ/hsqUBUIWSinKM30kUGRgOwM/SK5ruxpS3i
i8b8VPz81ymOXubYbTcTRNlYmZopBejOQJOaS1Yr9BIlDht0ptTZ6TgGABWFdxymqZwdMaYQrFky
8uSFNsEZZWVaABBzctXQmPGPaG3WJNtjP3u2GwUxaMMIDJua9xR6ezOFzaY/gO0gcf4tV5tN13L9
Lhxmj4Pt1H/1qBBC08d4EDt5Pb6rrWcarQ8azsHMBeaYyNQF60ZEA5QOWJz0e8jUBbGtAP9MldSU
KZ4GHZ+b8TG+NduUO+UZhTEBDCy8LeSw3j4rt46ePp2IPZ6D71W9f+2l7vTS65z1yA3n1qS5+B8t
nHHsHUyWZRUOQYKdFctcZfPWu7aWAaWj6crHVU7baOVv9B/4vu3Vr4J+4cgPdvBQsv4KR+jJ4ydR
Wx0ob0n7CX9kwiwiTloCfGSe/5/eofPU+qtOl/rbOmEKTXW9Ww2QN36y9KunF8+l4wn8tzVJFlnW
bh9X9eY+rJv/97Xew7kFhy8XHy9ZMxk7TR/QLHjTCFhhvtv+JLOu78dT8WZKPQ33xV48mPSwkzdr
m+PxDO+zk8qMXoUAc48I36czJgk8skxZ2K0I8GP90LB2H21Mpd9C3JdceQKFDD+XNQeVBvlg/k1u
hvxLOGtwFMr26mkhPiroHZSjAlIaLqjJ7UM2IQu+bYWVy1eyRv5RXFhKkatmZin/QS0Mm1F6NZi8
gQchnWxIrU8+IMAni2vEtV1gH9UyjeWyf6EfyLpzkxQ98vgdTGKE4IiEZXd38jJThfgxIkKtHNmq
NGq5KZbc6yhU+mKezRmJHhJZqnA+9cV6DRQ/0BbJDEhEPL9q8XGTIqQ4dODs705sdQEFl80Rw5DS
evRef+BCFUd7MCkk9O5/WRzYlyPTu+e940xCFk4FKHQs8PGZ90hl3sSVhShECW546GawdoyQrYH/
lVQa/LheDUYIiWGAY68v9IVPXv21MwaBiPyGUGK7kXjhNJn6XD3kMYph7Nb+zAdUAIN2AV2+Q5MF
0CuHd+sZlC/U+9rd2hVwg1yeqYLxSPfhqso2aXiVAVMatipFJkTsLn+iAfrupJ54OByf8kByX/wl
C3EDFieQwGaPguw+hl1uZEr0GvwD8yAp9il1Uh/efjswIegskXQPvvc7vCfeg2oREHNNgUbGNn1+
LnhwQKWOPDoz3zvw2MAdknFCHZfs3anMx2kh0qpqYS6+uq7ZTxgpFFAx4jlFXVA17hu6wZ+KLM/L
PrVY6A16gzuDP2QZ166VeiPCJaym41BFBAkMPmXZLn2XLWFow5zjSOnbwjJn1uGXoj6PLOUxoz2z
iYokHWq6eIWNhzRNS1iShoiVwJs8X3qSUlDfqa59dYxf870d0Xwk0f0nhBDkQx7kp+47TxdlhZCK
fM8zVUIb39fDhXrHie4X1EMJFv2/KftOUw2TqJdaDoZFSQTBrpjnAtjqjVVvXsRq3sPw8ZW9h1Vi
4rcuIfzvfAZaSiF1TRVYvkj5jXyFl2SVGSAAoJOlRHe27S+lOJXK7Sfv2liyl3fXAfBucXiwCDFV
uXRlDsY/E4uH+RWQoPv58S0/SwJzNQ9eJNNXoQbYj7GEaaSgDApExTrOk6LbJWwW4OJ3niSQmQ0d
8gDDRDWM/QeT1GYPkAlSjW98IfihMl/lYnfDY5mf8z0au4ehW9I++QCVYF1+4a3fIgcOfrpzN8Tk
UBqbViJveio+H5BFJ/5Gj5AgiJ7BWautCjiD+CoN0QzblA7IRRRxHE/fH45jMDEsHghPBHEdvAig
gHnW1DyPLOWr6oHsoPI2wasQfHRNDe0NGCevyHQRDJ1r96QylWz/mYfywzo17aQiy44vRFyyQNXt
YIVrs8xJDPeyNnpWPbPqW1WXENc13blSuMvgCuAA6sKTTWYgQzy5v5RTZ1o5i1kd/bj3Nwy6+dhL
UQ2yDLHoV1SRjRB3D36GTYwlyZDxH11Jqa5zGnyENGjeZGGQJK1jV8ptGB+4wFqtKbnc18lSmoov
+4s6kQrL+o77jRrv8fkwEy5Moz5J+GK13RfXlHT152rrsE4MuPoID4pK6OvjHNymhjtTw/ARLSa7
T8ViqjYpvTUmQl83O/QDsMZ7Pwf4lQI6+kIC4VAyXugUnECsrQzDVbqkcPrX1L/4uRLTCJDkBURp
OPwSMei7VfGvHLPhIxeWz+e9Jj5UJ4twsBjRmGOOY7dbKGoOvFH//WoWvXgl/HdieagTt7NE2YyI
2jlUE7utREm3VYFU3+/J7T74KGVE/zGEPL2A11BferBoNBpJ40xGlVY3tXFidgU2zduPOGfqUsts
umNNt5xLw1vDcLRfSLSvCj3eLp1X0ykvnKERY4z8zo2imiAZlNGU/8fQwxwWTU7Xy6x5rP5qhHQ1
354PVSu0Wa7ltqvi1bvnnKceA6gadmEj/wGnrH2Y+CGhQzZuWyam/pzvJGI4CXZojFCvvU1bbdLE
bhv3HhvAz5QT88kGYaZyH5X39VJiZYxmhdDD2W9CcQ3yN8NaGnWp6rNEmvsSZlYEXLHS8hnpDfW8
3bvNAJc3SznLydCGJPY3S1bBSpMo5Iii2korUueZBfRXHlazT5M2CQIjaboWRmbfLBKiUYvXf/ll
HAd/o9WPPzpLPilIo+1p05Am/9TwdUb0lt+QxhFAm9F/dsCY6pcdefoVoF+UrrbCfKKXCHW5Fx8v
fy9pqrJZYr4fhI2vKh9kuMAUGCBimq9KAwMf2Ul5qg8a6mrn0zl+AWriIiy2PkOO80xuzBuc6yxM
pWWKCRyKH+xiVjGTXljxIjEVeQ2vZ6/nP7hfO0bLk3Gk4Q16byrlHYEly3guulDAchHfgnTf19Jv
JNh6UjW3GLDd9y1RR0UfsC9l1+1DFJdKdMu7vOuKf0CgJZhGmkZ7Cvwght1M+iZZT1MM4c/3CfyY
9hO2s6nzAHC38G3RhDZLmxiKATESZh1LVWpNC1gF4XVMTMXPSIa/8JouZsrRoJtPfafb4movc38u
gKp1KZD5XFQtViMjDq1C2ieun0zYluMyeGmkggEF7zNvxt5xL4gU0diI7W5AV8/ECsK4oqtm7xHQ
6d6OT9ouSYk2ZlgDtMZvO35hHO4pK8koKp1QuDBam8H9P4qL43mE17xHGXPLuJtXph6FuKYzNd4e
EHobVtkcO0RWX5TQb8WU3Y4M9HldmP0J9vb4DVoici4cqtxeZ5dzVwmu06UQWfXcNyk4v+gY6F5L
dMGg7r4TnZmtz0a1QU681+1DSt9NzFGKNZ3W8PCeeFyjRQZnMdpC5oNYOjYNINRSDMpO5GaDry1l
I1cqAhmB4nw1MkcG/DXbIZMEhJo4VYDJeCZ7dGydUekW+BSrtHXDCF2dzTua+MGlkixgNv5WNhE4
sUG3FCFkdWMkmTgdvn+7jZJVyzLs6t/YrYcEaFhH+4t9tEOy3KT5GpL7d/qvLaa1gnDGAVgmvyBs
r2xUucAOLbM70RxqkcXtxaNlCba2xgpMSPMdYRDchaXaalUALPa14Ei4rZy8Vz9yur7YVMa34EQJ
EgF6Dc+/hq9Gxv/oHR+ulWHs2/+lusXgbJB1ZJtOkzvBWI90E1RWZTDQ3i+I5v0Eq9hjnRMLUcOC
xrW1JZJ8YMDn1qzZGaN8SYUFll09XKfoFYKvrSg/hvuklzvW54oOJquvbFi7xRkS/UDks3asgk98
CBxQXl3e6Qcb4d739Pb0kem61lDNdfBDESGrVaPWe3+qbCIZ3EZgzNcq6w5Y8bFfFaf1I6XwSOyj
7XcwNYiT/YBHPqyUH9ZMF1hj7zBMXqvHOSkeDyRmCtR+226M8FiNi3HJyQW+aij1T/Kgq9rMcfJT
95MnizVVvtk2MLxhG7ibnmux/KSf92N0CiQo+Bqrqjvwm8baDzMuMN0geoocWgLTJ+2gSpPMqPts
Abtm3o4PS0YSneKSpYeIOsa7qHIdbEdbKkB+5FbdsekAv9ayGV3WkhHjgzmFUG4WKUB1ubas+WMe
JVsn+JDuI4wkZRgWsJESKg71DxHhK8A7Yalifa8Y+PN27EyUB5TW0uV1B3bfsyqCqJdptoJlmgoj
xFipXPS7eXZeTvyC9LTDGQ+cYhZLqi4OeJp+27osN08jlViaOu07FapQk1g6/eGKSA/7zwnrcTgH
w6Dxq4beEXYpnmZcZTd+rMPb4Z8GK0oIrsKo6vd1MORvZls5K8YEZhMwX3hpuZpL9qXPKrb5e8M7
YHFRDxfFSFgHBnKNVJo93A2yf9xFRYazMUcO+B0U9WP9TBcbQhtG3NGA1LejQDkIX/udNleZerRt
zVafIN2HeZcpZqevtH1flBaP8HqfqXy32BlfJVR3Yrc74VYWE8IKjEQvqVr0xG0wa2LZKCwKsUFj
Hrlr7fBMBN47K4ON3LXukHtC3ORQbUfnbX6fcNPwVHgjmvNnoy82xwHjSpuHnO1LtoXxm8+u+14j
TqDk2MLykDONVmaC2vJb0/vUPvmgjeyIB8txVM8Ka4s0UceM5SGFyHp/q2fDHqQPhhvvWgS0N9MF
8BBEF0IHIgSwgOdXIOCVjq7LNpUnOBRyTd3bneGgPhU7Eb0FV/jrrADm+RiEw08qPMLC9jx1UU9J
QpFz8N46PHLztN7tzfGqEgKJ0dKiYzc+5d396A5kSCCYcHUNyMPyMDB7XFXBtEN90ekG/QudEHow
EakXdZWuP2E8/zYmNWQQSJfrGM8+YqgQmepyq5HNIu/gfPX5bCDIP2/DKuzcZK/WoyQ/VPOlE2RF
tF32BvuIY6d2/jIVlm7/w1d+ZreFHoSiCm+sr9XFn5gDDEGg+WiwpE8WSXitjs6/qusuoCnZha7u
YKITl9WlOaoYpcBVzskI21dLyNn0rbu3708EMHKCR9ty+U9XhfvPo9vvQn/Rc6siLAQlgpMaGzr/
Eul0ueAef62Sc7txJQpp/NcCUxVFi4HlCWBRRWY5JctAlszNtDdBt7Kya2klyXnYYfoFG7lZngGz
aiGGUxiesYu3jJ18DGmv+CKH1kTYd9ppmdfd9Xu1Minq8GQjuQifJAgIDC1O7rbgiXhBl9FG6VLS
dbQL5Nsq3m3lQ69VywW5/5kbqIXmt+uFFTYSReFyKxAisRhzvFRpqB/hK8GPySdCUxHWGJ6kf8S8
VO0pCXCgpPXSTilxZ4fY5tGlwaepCobIO/O/ILqd7H9j8ucoCsqvCWJEW0YYtdtbK1rgMud2ex9+
TF3UcVKSIo6K4LHbz9P/i8XGy/+J9JUgEiEFGdfHLTQu5Fu4xH+3VX4yoa0aaxHJWCge8o8kCS4d
XbL6tnmR1srwY6yca9G6UA0FNiaqb6iQ542lYzFl1rKkufaooCL4oI627fPIu1T5bON4CFdbUES3
VbBLKHw0nVk2eJHewWIuHSWm+EL2pGpkvS/rIfRfQTen7RN6gYlYgVmB8BV6tyKAFvSqOT9CloUx
MzeGboqJLBC7KQ6wmX5WQydMfMWwRp3Xc5357E00Ep2LttP3UUhgucoAnMN6Y2JNtNRKurBfYna0
muNV5dhJpUW5ZW4WeTTHQBTK/Z7ZgUgtzYCfScDuJVJ34f2mULLebR+K0xMQ/za6SfneL0oW5yPV
7TVlsCfO0g0MlANOXdZW5VMMqSiWvb1SWNrFtxYSnwvE4wFb6+mlCRItZVQbzkmVYXJhdBn2+cOd
8LUEklRcFNqnZolCWlzXGJuFhQ1hmVKX9OrtSt2sNpnywjdy1tiXed14uUxTv2cWWTaw+NZa3xTZ
99VZktXBoPOiMG5M/9cDeCrNMgShhlZhZOkoosz9zan3QEB/dV5ZaPZgUZIeYyk+UKEXRd3X3jjS
Qal0w5L/tdFPdMn9Uqkq9zhP8DLMT5yXvSmkY//P2cGarkqQcFp83L1On5S9bylZMgZMZPmcOOIM
OYa0uVcK+FFVfBElFYgwep0ivCGtB8yTazYIZow8zYPDZSK933MKjWgLCAK/VI+WYMGvGRt9M3Bs
Xot5uPR8DcjhUz0pJEEHNe5kuOMTVoQe5khLjIyIQZnKXUERUNH/lxPATxbCyKQO37HlASQ1NE2p
2K29x6nyeh/gM71kkmHc7pVi4nFCgfXPLFL7PwBl0GySF0l6KVVw3aEyLK+dIrA2C52bFTHwPR1P
MKdEJ95vKGJuY5ZepqIeM1XVAdeUfZ/YOvh3nW+RY0iKT+HWL1QQuVrzJroduxhrRmt1hD4Rtep6
wMiMbrpI8STjq1ZYYofOSY192RxjXps1fOcmRVK7a8NnF5i/z1mF2cHwK/w/d9q2buEjLNfkxKYG
oulvZk4Y5v3vzDX3Qqm6ndrNqfOEzP0M3RcRKtybECOk36SQl+RIdeRbirO/t+ckVlx907pzNzm/
/JhhX2NPUkNhVsNO4r0Tr/LqLKCItgSZtS2CZVGsLHpTAQBrH671GxhzYhyuhmVmO/WpdFLU1PNp
//0/QWV0aj7lyZElKD6yTyuI1d8TYyL6JjpbOLngWAC8J5ieZImm+f6Qh0Uzy8Pj/CFIgqZ3yeSn
bGDvLzflESHXKCiNCykyXae2I3obo9jxf+pstU8MGANUcDUmt2JsCMJpED9hAe8/6kz6sMqDXTKH
ShdoOjTHJSp+RXFl9JLYnRRZH7VMBt1BjwS+XKWKpjGQgOTkKHB/wofM2V7AAMkn+HPEfDCgAGW+
1HDhl2kt0wg32iT41PnXS/T1y5rHkUFaJ6QXiVPEweSZ6sB3IJrayHwXaWisxwSEJJOHVkwxNU4D
SEQqWUVsQnSAB7Dfd+aW5rkDL6eLfDzWpkQlwkWVzozawp7PiU3XViD0nFvyHHaTipXJ8wcIB7Da
4l0vWmsZW2TTl/JrlkM51F3HVFYzjR1ygCw7P2AkaxQno2M96NqWlEQ7kodsrGcNEtOzPj3OC6z6
hNQuwq0f8AyM6WPkqNUIsbE/u/s1W2n4x1Cgr7f+AnJl7Si5X0PD1P8E4xKRj+G8+yfDdDp45VfE
EzYbnBHpeWmsYfl4o0isFVVb5GtmrBOF8cjsH1vQwzZDAvBq17xB9f3WwyOigdy9V3AncQp/ckhm
PENU/NUarTaT41p1kRW+HRywMpBtEFaF2u4MhhX+J1k3G0as34zkQ8tCvc+f/vJt7dOKanuECX4U
fKzXEGmCLikFXRWiEHQLi1ZrZkrSQtHClAMfh+JM3I9Zt0+5piPYpgyU0wxuWDu/rOfjHY4eOY9M
J1n/JsX3UF0MAKqj8yoFTM6mEYS8I1HNrdPzAlhyPdV7yYGNkZWyRWWG0g2f7281kK2yAWLovTcj
8dBYU69OCBRR7eDnxPhk8dqAj0vgZCvmuNs7gy3sF2x+22tLfNGeiLimTuFCCa6wDC8mtwwZN9Em
YsL+swRO6OgJFdgs/xjgeyLwWISec+xjXwaCN4I/D6kgUYpaGbA57ocLZPFw2GqlQzsWJs76qBn1
I1Ms33PphvcUmjz93DGyOFLboDG9JmFKSBUhOdmDPw1ZWMasZp2Jg4mZiIl6RLoB1GRjXZbd1B3U
d8uXCPLlvx+Lsnxq0sFbipGIYthVtRWCrCXuMEGqfvI7MCCLqaCcP8rGtpsMYblR2jwN6C6ptbNr
fI0Q1JaIBwVvBrJdfhDGGMQu2dP16oEaxbWu2dvDeJqYtDSGEDZzsqw3AdQIV0hVMh79/++ksrBb
/l0Zqw+dTqdRfdGYLu8il2Mwh4x5953ulSjo6IOniFScDzw+5PwkWxH4fARhBf9oHzqcSB53Spl/
6JPwWECf/j4709DjHHn1GFfsFST7R4tkoTNlGak1tSxHcoM3STAXC71yViDDVzPn0ZFgdQO8rEuc
qxl0V+BuIDetJgJ21eAp1HBEejdsMrZz4NdELyb0Frvs8IDwCz36Trnr5yqv1hnwmRLizCenzD32
mYdfsflzYJhqNWdXy6YwfCoQFA5IqzMnW1VG7M64RQ88Z3HjoLLf5+P6e7dDxvWFCN1S//JEFHcH
t4nPg8TdXeTShme536lrcOC/Y3WSruXbADVlmB2Ju7EwH9kWudfgDWudwlCzWfUx9Y8HgyJo49Vo
qh+uuWVZqZCU8Rjyt3qFfO4sa8827aDi3zSdq+oxD3GzYnpOaxmMV6mNRp76beiEYR5j7UQc5R6v
daXcFSCKeD6ZlVyiZjJIV5y0GsGJHYnGwrFJIqfH4N8cWNjN52kj8Tn7S7N3z079b7GyMBg6DSfO
gvbmMmyQ4saWNiNO0+UplrNgm351r8WZJwc5wM01F3prhgnopbN9VsbIa2uE4gqk4ipLbGOOBX17
IZ1e2hVwdkzOktoNPudaD5dvrr6hDQipZS4Vh/olnaT86gmawKRWTypXva+aYG34zwlCzfCJt4PA
zYudgU4wkdH2kVBJUb7YbqbwrewokSGJ3uaCKYPh1mnUMTSpPPzvWaYLDRREv1VivJrN2rcAM5Ah
oEG+9Ay/lISC9fR+yH+tWJ8WlVQOMK78DpNBlKXMsa2hLD5rqSJUcAawkzrXB2h8w8/BnLeWCSbm
uBgz3bjARSX9maKmQN9qeJMwpQS+SEYTgYsqm0ZUiOjl+RRrDDImy/Hy/cAyXsRGmif0azp5iqKX
5+yPLM1mJ6RhGwFR9v9NgqFU2uXmaMfYeUvCOzY1ZCzbMOZlgg97m8nMjiPKLsLaSx0TRga8PmYF
d+w/ueMqm1l+QxS5uBtCMQMH4xH5Zptnf+DvEuoNcV80ISaqInitztjeQwMJhSbsJWmmd68Us9wh
SHHb/z45RpE3d2kBMverQcNxEkhxrpipHxKJsOirkpuC/bf9G/8CafS6gHTbJuDRoJqerTWJh3wS
auQfSQI7atcQYVKIr6uPLnDn83hY1up5ZKGY9pOZ0KetpD1m6PBy8ww5J+GR30KkWoGC9uWSYCax
ak9ZEfShaAb+Z5/2SD89G2EzXY8o4xjzNfNO8pCucurZll9d4gripaicbu0u2L2BsE8Tqrzg/XXg
LZZ6Po9VTMmWjd4DBR83rQLFycwbCP9nfy1iztfN7Vt3dg90w6dg8MuCc1ZPNJJTj5xI1Mt42OiE
Uj71f0XoyaaL/X4h/4V5Pph/XxrDKgVL9gz7ChOpooOzybDgCvd0mQZbgz9e0+JRWMdEwTAjfs7Y
Asr/So3GTn5zKXVrHfdBVZ9D4ZD1BZtb4BF2h6BIckTYnfh5pKEaR6Mu639A0I31aqR4fwJeL2NW
kG42RhVcY4PC/X19A0zh8zyOxcMqmthI3WLbQryvVNEWCsnorvGXSNXxsTCy4mqRjZf+dnWEd5aj
WZD/ZV1GajF2NToPBc/dEy7DaQT++UWQ5RGn6UhvSCSLFbrVwYykLsklxOZZgKnm2ZPruBGixeux
oQVlZPnRNfW81BDD6U1/lICpcm5okOVXc3f1ByG8oMmXZ3evkvzrafomJCn4kt3/j9kVLKIFlhml
8o/jczyVZCER3IHsFzTuCIU3PDDjQGd83adt4QemRCm3s6FL9sazhVGxMo4oh+sFLqYIN+DvJABe
olOTyQ/iZTZ7CtUMv3eoG+Uk2pzXsjEy855E34e0wucKU5JxvjGLRH3E+VzPBnhtSACGmACseEaM
jc+Xyl19RtWtuAS1kSWnIXqfVvxWtK6DkD9BLHseGBzqBo5ZNGAwui8rywZ1pOeP+UPmjnYuo463
gjpBjnKiG1GsV9ihUmK1OoF98AqwZUbk66m10nDdkMp0tDOqwDx2UEVfxqbOP1tv1yzIrd/3NQ8B
mIHW4plOhcFq2cjDlZj/RC6WRwWp6wr4Due6MJRWAgb4Jt0gUpzgL2/0W5tym3/qzHPiW829zxTn
4Ud+wFvRc3J522LSmGHvQFfEu93IFIVndBWtMHsph55y92IDr/a+K9JIHDXX5xPxtm+DBFy2fPUs
utGcsWtE3Fs7JqhbEJ4jdwSBvWWnvGf+Ba56qfzNZ1RVZUSpuT3YV8rsCHC6lvSoTt68w0+We0pD
ZFQDw+1tSg4veOXH+UxamSfmHELYojiNn28w9Xdr29RBfnr+sNHKcNwmTugE8R97P6iGbU+1rgCS
JYJEo87i9FpvrDwL1jRfakw3KvGGGi5hoNPwUpmswB5ouBUHcCPg7AgtyIiZ/CrXE8KlW810Clwq
zdlPFNcXN9UlzRitnO8BuCXYRkCiodYhUngKhi3Y4NBvvQPd2UgfRcwuaqxEcIwWK5TBZFvXhN4U
XN0N2SneP108QaxT7C8tN/KsDsL+1+YaJFF4fo+C4+xH69TK3r9ij5WYTKj4sNtmBvWi79z/W4Hz
uXI8/pe9TUEMqVbKEA/itlTYk3Qp4mWxqLNHxf+2fNFXMn4bdrghN6jfYMbXznoV+Uj1pgs1rgnr
FSluwSH6+IKn09GM27jQeFgl/cyIgU3MLsiBIOuli7AOxCLepbywIj8+ovZxLqzqmMd/xMlyhW+O
jtZGgJJzDKD8WILL827fVjCSr8R99DqEsWS9p0QbxqjNLhb1LL8jGcjk2mfZi3dvMbv79shkSuMt
N//tACzTx8+ObbkfJi1Kz85sVI6PX0eMsQpIAXLC9OdXtYmAm+j8h6DGMF9LoY8Cw3KRkxEuC4qw
rh9U4OGAr59+MjB4fkz9Pv6yGooS+Yp69fX/Ivu+xCINaR7lqUxvAdQ4MQlOEDKsxksh3mEjKkCR
pxyf/fPpjYLSJAap1ptA3kKTkphCk2FJGN6nPqKtOSc3ByFy9bQhyFF56DBRhiVxeGfJotHnfKcy
rtXpVQfpFvvDZzSaSKvZvPLCVsO8e16no5NMHdHMP5INQigDgMwcfJE57jX1JUwsoNw80Zmvn05S
6xrTSitFAk3r8utFUzfSqa+pn+ur9hDEQGma+ZqETd/KBOOzA90acMY3tDms2XfSOi7hp4XIHHlS
uwicOD0qq+M6h2z/fSJxK6j5RtLCyYthuHt6nbtiK6FlqAnE5qw6fbW72Zx70tkHDQqWkJn6JUAm
ezbXDPTJhx45xIXGoYoZxRfhtc60TrmqwU/vPczN4R/LUol4ScSKCA4c/Lh8nnm0t4E5qOlSWtgJ
mSmTiaoAfguUY6SWllLflAMWWQEgXeeGaabqroWr4QB/oTJAK5S2flAtRqdZTmgoPrQeiznV7P23
BYH//1PiuZ+NcdCFMV1Ql2dt20B1YQa263JryFHxAvgcvaAnNFB4SVPm+SaVByoQ6jpRqxtNzoYZ
WRjghW15OJzn2qi40p7AV0ffsp22SQ9ACGYOyZhHw4iq8U3VSREeRquug3s+IlkZhzfBYMcNavy3
bazPH89cizijuCQ5n+htskVJ7F9iU6E+z1Ex2V6wqcJQkkSKhwuYSGcRcOUiMvJ1D1yVKpvUHlSy
iyBgqX4pykU7uOIENtckqG76p03kcoEPRBRxo6yc0egi+H54vgL4PxDBWLLMOStIlR9u3O1+tlqY
tGayJiJURfMamICVYThO1Q8q1mqG66K9UEzVdGWY49FUcbS5zayOBbBFSB/BiKtuO9gqI2PbPTUX
yxqEJVmxaPiUAO2yiU1f+DI1pPP6ksysl3eADg21h4T0kxWYrIQkXAhuJpRgYWGUVnaTM0VwBccf
gIWCUZbjT6VgTMjv59HN0K3hgMkgFSA2e6NgEF/n+xxVwBjZKQL09zPAE4e4CPWHZmCimkzMT1oc
JGquLm8NqS+JL9poUr8pMpWEGO1wjru1tCJA11yTq+qAext+Tp531ZTa1OVtOpMeKJKLidjUGM3/
FUHYlvV6ql5HIOLeZuFkUgg1ynQEqOc7orDuG1s1lbKmS62+EVg2nkTpKz/caZJzw4tKB4cNL8Az
GL/qfHTFYZSnpiCwKQg65VW8ohHpDl7LWBbLfpK7ZN/OnlEOb/YvKCl0T3vKAd+QVnBI54RRCwX8
dGitmz5kXEbPbVItaAIawYdfIZe2JydhhYSOnsEkGErvyi2EZqmmVCw4ygLd8Fp9m3vbt67buxiC
etxUqkHQlbTx6CHZkPrQ1bt/TC4/yXsu/WmYoTDuGhbsb7auXjlwoUol+2ttZzZPJCSsXBxM47kH
4SFosqwqMA6D+yiVHrDEWea0TdjdG7Aydo6GrMS7QJzb46yK2oIUlbEd/mW1Dd819eB7rDA/UvJP
XVjjv5HRPY0gjM4ETAuLclrXxa9iHYizhS1z48pPxKa9GK3AzVxqF6b4v0Ax/6zUq1KxlQVsIqsn
4D6GcWWCabOb7Nl5vciR/Hjt4ue22JcVZjIdTLm0PJmlQq9jXxKKYB2aSsArsb8NUUy8zp9TV5eF
86Yg6rJmNVARVyTGwbVvWOdfBBo4aygXhXNLRMpzF2GbrbZPVFwY2Kc94AdEQpn9cFqIGBbFmWMg
TgE8DbIKNdjM+WWW0+T23bs/KGqYcCusdsWkNmFGaQX6YzBtIGIGEfxGnJVuWhzfyMRtW3X+s5pp
b+9/lBchzKMsyNcoHp6DqkBUq4K1bbSZkgd2FXoFsLNfJNhho8Ywx9eCR5klRLsIGvFQ7Gcn6fd/
5Bv6qP7rgoZdciGYcFLCu3Fmh5O6R4tvKZXXuAI5PhTScieED6RAmMgnEN79/dd2itF01+4aReaJ
tNnCazyommI60ZM4m68Zi8b3l3wUVZlF7u/kJiih11lUjDOMbQSWA1GMdUT6UDeNoFlC9zDSuuWp
sB+QiWkDiQB8k4MjK5N0GlYnEx1Y1dfxYhPOUDdJh1z2P9Hk7itXOjbngB4ww/3bmmuRMDV+2nkq
Ld2jr1dCuE5k5bxLEq2SMj29lQ7fP1/vM1ubrdtZhsx4t01e2ehNrN2n8rVXbTPfCoh3mFsSZfVm
vgg3YA9P6Kd/jXV7CGb1nA0YKZxxSqcnrcmQIJ1YPx3wLo/eFynG2Z43Zw1FvnXaJmB+gyvRNnhS
w33k7KRQHENykjaYFb1vLOs9Y3CLRMGRy1uIaolqoCJWauoDHfJZnMN2EUbanaZ4L4AEURCKRmeb
aizYgBDajJMViHyyzbrf722V80RdEDNlVkI8dRHk4nfXRmyBPzAtNyxny8CeEIG9BU70QD3j/98g
72alLOwDFDpVZpFOeycl33cVeuIXG9RIyVzngR/3xAmlXyDt38GI0SOB9iEtrV7mBM2NncwV33f0
zUSIjF91ERGUV3tSG9WPOoRCkf2OZOouVs4DtlIDKhYgaLg9c6MpPRJwR1QX9UNdM29ELyhFuuoF
FMuhj7N0y90H3WMvOrQDwfvDkzTNmTpVJt+EnyVZyIs/nWLQ2ekDPq3MinhTCQKlsCNDSF9vTyr5
CP3g/VPY5yrk7G2qlNJNmhj2zBDGx4vxpKty930vK2HSpMD3ssocJUU4JM++EcLCWbYCdih4b4c6
RhvOmbdota925atXL0mocK0ky1yal3b105tQOAX8aFp0j8d5VqeobsmBToXzBYycp3lFkI6y8oGx
/aYL6hrG5l7C7zdRK97pJTupdjp9bCLDzUuUJqAsntoPEct2oYteiicHrT5LABrU13bY4n0paYkd
L4pGx4Ns0z9YPiRtm4tdri6+LXJzmw1YyJXjv4SYiQTTxYM+AVFQq0/ZnBgz83lEn2xrnlwTXK4N
/XHTBq7vRMf7xeViNX5feFDWQt8r+eUpMatQ5u4E2LHgELrdhTg3hE571O2ImPeW9n3Ev/Hh7ZJX
WOS2xhtxj68QjyGQBXTPQ5Ck6FIhs99Gfvus5b3dBKAGO5/K8yuJVzabdAExg5CxkrwePlzl0dmX
E4PJzmN9a2+4Lb2FP3Vm24dvvwIIpgnIjt+Ynlj3p2oBR5aXWayZwJs6QIFJdtGMNOV8fC5GDRj6
LgEuyEfOMQr51fANXJPtwJglGYFRklUiAcYzJRb8Wxja10qo3HVaFs9O/HxRCesCTRC6U6PBAl7p
oPYCjcH2t0IZw6g/T4T6TMhlfsNjHjsuJ0Gwt0ot2kM1IQhgRXh1ntF1S81G88r5OaHtWm36SeK1
BY/gwqXpLKVtKm029BXqMmHjr3pvHMk6Z7Uo4zfkuS08bB+bJddfJS3pDqYhYpiUmIl3hPW06+ML
qyoHzce9tVlabpuOU/47XquHwNKzSaHT+99XPJT2qAJoengVJgkVZNDMq6ysuklNTpxfmGYCTkeA
6Ba7yVYUBD4Lx0C8p0/N83UtCImzo00hlVzGAhOGqDIjlsMV0REfGAh0D4qCx3xrAnp7L91rsj0U
3LZRUlDS3zv+RJBzwqHfjM8eN7nadCqMlgNfpqytdGwSePWeLkyfS/JFaZbctlqzoO05C5tdH3Vq
bxEan8CgM0Y366qWpu/cCEEXx0S0j9kbDQNtlHW5EwveHd95kCYHAmgHt3jXUEelu0T7mZ3Hn076
DNUWbIb0lGSxInOURebru4GDPmP0AHprPQxiWJnMqpDISyjDcqe6LvWIAD+WdQVq2X220byaEQuq
1TW/4sA8N6zRgEu/QEck7cEockeiPISVKP4l7WZCrNkfaVC+iAiDMxEoxFi0XLoQ2AMc8g9/HbzA
hHOvJN2sfSREdhr2AzsVNl+cPFSXLWRRgSqSvf0t/HKGen919WgQXpUtL54f91Qz0wfVumOSdCGj
FmOr11SpmiD6JckG9zn1uewECOWLDmAjuknwmf/YP2iAXCCp25yFhi+/6VkQP9pgXoKPPxQY+898
BWx7T741je2mnY1O/FUHHrTlFKGvPcyd9f+Fjx2Tl35Iq4+1b9YLoCP0YPbhxQA7q+25bpheDtlG
g3Ze80HoSGghNunxVm/VGYHatRS98yBm2bsyBlctAfzvgXBieO30vuysRMPG5/FNgICxEfAcRJ26
cGLwUaLc/BfpxNWV+XY4KTM3A7nwBEu+RLqxw3eNkrzuDe7HqvA/c+ZoATq9i6V5Zdw4qN8vJEW5
+qZcjMeV80+cVcZHsdoDj1mJkAuqbBmmLZfFuiFWqUTR6sQH21eKpFUVbsgq0WXivBDw5/L0EpC+
PmtptvQYxthZKlT+xwaRMH+8rIfAE9M4bpZTZ3Yz4RM7ehhsZ5lei4jz18nzRmUvIFMEFFMnaela
CB5vMCApEcXWTp9B518N+MBGxdvcQfeS71JdiFeMHe3E6GImRQRyoRIyVx5zR2SxrmFQ3y6vVPP7
0Sg3YaEiysdZSKGhc8+7/vng1XoW1OEl3sK8TdBmVnKRWuNiKT7HLHwZQXw8jTgRjw81DJlp5tjz
BCaN27O5JfQ/tbiMjTM9vjaGIum6+tz3y9SHqAvfe3eyUyrknqPE11dydPZ2Gw47iVsEPilN9b7e
727syhal8dWPIIKMc3v1x6zw9+umc5Dt9PERS2lYupacSUp6Gt/o4OMkEEDSA16TBBxBdr900Un6
Vf2hze7IA9us8iHouHxAAeWuLWU1oKm6pzKGfpTMRPOS3e593s/iMQhn1EydZjZp7DfU8kU+PCeQ
+1Exw1xydnnUz0HHITaqcqtF9xefan7OBNqDLj+zU4AErq39/Augnxcvsev7MwGK+GcpoNSl2VRK
KS1VmSLY2RBb5LeiQdQl3ZCVKwPOOb70qNN/rXN0xxJK6BRqhMTOLLXIXwM8cPA9161aZGShMgmk
vrZsT6cskxIm6/IB0EYn2SdrB9ElnUYvBgqzulou4waaPBXoLxM2qfwtox/NCbTq+yYHRktZCLb5
mce2/StmINBLsk4SJmbH52d7NlH8BYB57gOLd2E51WXvB3HMVfB5b2wiM+rZc5YPoyERS8FHQRvx
8xI1rxFemx2WiB2CV6j7lu/R5nb1czjBjttgDnXuYNyq30voCDR4+Xc1oZKZHHgzv/1v6mDE/VxS
KiVUCPcvFYWWEqt36j0XEuIUhHxJl0kK4nzMrGqGgPObVI/uZgbJpszSTOTRiwXCvfhCdU0E0Mzw
HAlTQQAwonc+IY7hFqggfvzqbH2BJkv6Uria8S1uMxhX+ePz5NfRhCAmWV6qu4g3km0OxyIQxxvG
KdjZR8DiR18CPwGznwcA5A9JhqXsJbrp/q+gS60NsrEJMy80FpRYDJGwxuYNgOOtb3kpy574jR9I
7Eo2TP58fA1XNKC0oMO7KvUcOXEZ82jFFApXbt8shSD11B4R/AK9A9WriidU9x3BG8wUYES7T5OA
Zunm0TR2Wdukh4hVNdJuC5xA5vXQ+Vt+jiA4AopAB5xc9rnIo1HkGh2xyYTMP4TwS0aUwWhrlMfy
8+FpEhLmZ3I7qOzyNzPetRqRT0ZbpoTusXjj7vJ2gHUmbPgP9yUIGYejiiWdCCWiJby16zeABE2N
K45Gum3FgCxfZWf9gm9Vkjd6WbzKMwEUYYFJPhMcEEA7kXjQz2JZkaZcDaLvOOx6rtXm82t4sa2G
4+ucqUon0+cx38id69t25dZTU/gJK4ycoqedrYi7WURA/iDyvWnovc/Wu0VQd1ztJRyr99mwoP24
u9xIbihx8jVsoEfMIiBTFeGmjWcOBuW1zRizbqhZFRGZ6QdU95g+8nZPlelazMfCQAKCaQgoNH8D
NDigXrEkDFJGLlnGDtgO1bJtJYKiXIzbOnPziJ/LvJC55iTDc8tVFBQzRO/P9UHBmyB4KzF6yeTQ
qfJdh/71TNIqnftGSqZzdsyAU6oJN4bgwpx2iV55+tOvdwYpgP5U+RMxunj8VE9luDfilZc/eYDF
JmMTu8wOpMiyYcJCOzrxvG63Fr3yE4UFdrLUFp2aqa0e2Pw1SBdm5OfFVh7vb29K2nOkAXKhxO20
FTPAk4lAl5pJqyRRB1jox0lLZHQIrIzrvOQSeJMB20r0KdqGH8tvPBY4sTYk4e2tkfOk7fb1AP3o
b3l7V/nPOeXYIOI1j8NJMms4Eoof7UjjlfMInkItOEeQr6ksgVYCv0Dq10blmYqn3LK6ARoMwvOz
m6SG6qyKBfkx0UcRbIqaAH+MUed2dBuJ6wRfdutEMtsqlTlecDg+N6xfVFYwqGlDd0q89vvnWkey
Tkv6TsRZjV4kQ2lyQBVCAW2SMwl8Ys5LCmTu7RUJqSxjhOkws3XMtYiUUG14UNmD2457VK9Gntwx
2RbvGsfa/TEKDfmpDRRwYm9dpGqNIYtfuR1nnLh8dmG/QfPa+NSqEfVdvfpn7ZITX7UFN5wspoYW
201IzgCYJ7ZlNX/uK9nPSB7dJ8iNTIoiXsyfKzi4lIWq4NcHUqJJtZUp4SkfLSybCIRXICUMh2pX
85CJOCbFJJXugQBgPme8ig67bHYwV99EmP+I78NJCN6uNb+r5nIAIn//wymuq/N8wovIDvc6OA00
jV1z3oVW6+EG1prLL2+fY8LG1JZZ2u/vGixs822IA7psLB36yBtg3HNuhw8Gct7DOGYSEHuYDT4P
oJbK2e2EDbkHSDdEBzP6HslTbPMiBNMbhrrYD7NbrzIX0MXRTylGKjeglZ1xVv6NL8GD06aFC8+a
NWqAFfa3qjBDQ67IkNicgVFon93+CvYGK2tSBxUw6BilhP83D7gxVZRJwVZYhOAO7Fhdm2ZKuDRz
AS2Ew+0GwfqHhNHopePvJXEd9TvEfNBGizvklVz+5XEGAyR1VQtF73m0nbz6s286tRkTTc0kvsUu
4RTPFPcZ+dvPZJryqB5bNY4iMzLObn5ugfXjsaJw2p1Vq0ZZT/KYPWU6QL65aM7lSxvNkNDADFVr
0IEAEVUJyRPI72AdCdM8Hh6aDgSdj7baLws2q559a6XQoOF23nbKDUStKdaHn+7zsXqLJgQOlhuh
BZUNCjx1dk8QD6hcNQu8XcAtmuoC+csaPOcayETtGLVWeMPvOc8+r91qOhPzVIW6KyZjKgla3hSI
ivZN92okY5C8j7n75wtIeaP1UfPMYn6Jds/X5qP2BU60Xw1vv6BTbaHvBHMCrZXEKtXrz7nLS3ze
yIk7FfWvWR628o0q3pR932CCdCcAGTDVlHDugnxrkWp6y0LJB9Ri+4MzFEJVZI1msyPWO//v/mN/
A8KT0pLNRVc3g8P2zxZffF+r3LeD67uE93c8l8A/jRb0Keb+xxVBLHjDbCCp5iLnOkrKOXAnWvTr
WnqylcUg5H6E9ttDdH4rMJXI8Ab1UaRbDOlz5wmxfu9Axtr1ZtNhBbQENpjq9Flqo/KHbm23xSBw
v+LUXl1C0KGuLEG47obfJyAE4QeiOM35pzKqhw1TdJzA0ovB8CMEBZsKOjq9C/N+gilNIjEmIc8j
TPX9kEh9SkOfxLc+AXeZKC2/ZVM/7H9LghAiT93Ah1kyfUzy+Uu58atAg+TsGJyArLWyX76EauB5
GoYGSOizZq77BbugnEskQNJhYPsneiG824K+watY9NWC3J9Dbt8kiPWk4N9oZlmBog9d9IrRAx2g
uSaD9CAxi4RJZ4+lDPK4vGgki1ToawOgggdI1jB+DUVbd/KEyW+lBMSa1ihVu8OXOiy1aeh+Bqcu
INghjACsZp0p6no98l11wnXPvmKakLFro+m8EDJCjk9dEQ6kUfpcEh2upUM+FFyabkJl7vaHZKn9
P5Q02muP3xj3YdCgx8UcqWcJ0ovfBbshZrlRCFhgqbaSJ0FX/Ra5DzI0rBrGsKyWZX+D302c7d2+
hR842EiJQr+pDDfpcWoTOqWSW4GJf9KaRvcenGdVgNntiWQCdYToKewr0vrDAWbEYfaLJd0o2ge1
Or2D6mWAW/s73blakTS51xhBdqcI7hc/WjN3m8ZX53ESDfG+lANSB3G3VYzeuAClNzMRh8uKoE87
+aTvFm7axnRaorKWWe35Cd0CrHeK2Jy3myWbnMSXG5/iDlV0j1pjQQt3rx3RyFvEJTn7g2/ERcOb
FHZolkj2RTyJ2psxsN/9FB/wJzVg351eyHA+jlhFa7RU17kpb+phZPlisewES13BEKHPVrmmq/LE
cAGtHBfEmXb85tc73Bs2cH8x00kxH6VoDimaCp11djnyDCdG1H0BeUTCxNPrk8YpJKOP3XL2KmqY
dSF1x2TK6g9CJ9o4wfdhRFzYTB49gD/mrKeqwyGzFII3jadE5esR7eT89eth5OpqkjDrCRmr77Bp
ZgoxkRangPQBznKp74h6FN35zcApMwM64UxVqr8EDaRG4UOt7sNntTbG3U10xm7y9pqiEF4X2wpY
6qHIiEVfVqHXkUiBxoUIAFnXFIIfwtumnvAhKr/hyN+4WLevZPrYTIRhLJK2+xBsPj9uydn528Hj
0O8yq0hD164OmpxTDHd0tUi/YJGlYg89aq5Zq11yYvF5PWUNt8wHodLM78svlZsLuR5N+uqVVfDi
uTmJ/Uwa+ucl99ByV9RjuafXsmLLPcZOiJttianttnHAp1PBgPd2bvQlDWGUyr621m+/9XvN8W9e
i/L73bu1RAFFgIcyHV7t0T/vIz1Cj9fTHDe23znFiJKypXItidGd+Djodv8I9US0CkCHstnmsLyt
iAQxWeTP2OwLpnRoAYX50rfpxyCRhqqSk/8BajA3mhI58goovd93x8xxGYS/WGGWijZY7JjS7Ftg
lqssUzdvCF5IHHsvthI6r57g8BmoU9ZhaWJZmQ20lpnp4ni88Sa+b8LU9PtGo7E/rLFCgFzYRB3Y
I7xl9p73FuNxoT/vMfuQCHVQp/UDHlK3WT4fiNo4ExwwOQoJaEhZxNduwIum9oyO+lqP5IsqZaSL
RCi9B4s0ANMLxOLaa5o2hdVJhQwftaZXIV9Q/O+sOHySaHgcN51+Yj/zbjS72SaNWyIgMxnVhQzK
E6eZMEgSbgu1dnM9OJWOww7lDD5ScYFyINLo0fbGhpb+9nLkZd69l7sz+FnOZTFVziXrsduMx3fm
c8sV2Zh+rI9O28zHnu6c8Zn1FPaNyjd8u2pyn+4aH6nAi7RCVvBbjudH0f693+U5O2yGnFJ9hCQO
0Ao6AGJPiiKKmjzWUiVgWgX1j5uhq+bAVziHaSwbq/eqNzLFcAYQXE8gVI15iHDCG4OpO7bjWn8Q
a4AmnjKGPaVBY0nJdKR6F870/dAcvP5HCvyy8PwNahX7QDIn5hgp98pBxN5UVfAChyZ27xVo6A+0
2xgBcb/qvrGqpOkUfUnR80uqw+JmaEN1WNPnl9Ua9Z4UHhyfyapqoNoPlNpyFrZCzMwGnTKfGnxW
7PKO2l/0AhyfX/x1kG6LnVolQpDe7usbWn26/IBGrdu15Mtw4QSqMzel2A8Pu70rWujUQfliSRe1
bPARe17QSRaGLHvityG4jpfg5vD87ctrsidluj961WvvsyHiiVaZQ+tvwJzH7sAPUxiiHlSaGqi3
m7PqfonQO3oUq0mdVSO1EX/N5cf6HHEQfZwIE++CYlDTrWnvb4xOgidoBB8DB+0g6a+TqyzfdTif
DlHvScIkBFXs1WXr6ZdBDWXIIV0NE1iEEJxSb06VwYoxIOYwvT4eHR6dSyRz9O0iFEoSrfOSB1nS
fxIApGioLc/HaqF93KShkWVDBv7qq5qT4l1SQFlXoAPTf/LCMZOo/N4qnDAxFfupGU8KZzIvxWYS
dqXpvuS+tjQ0k9p6EzvWUble7BVcDKo+7SD53cTgUNVjw0Xf28goWTq6tu6FmjgCpKjQ2jt4pATw
nxxz7FrCd/gkAE25azp+TAeF07mkziGPHw3V4xP6lC+0WB7kvnPN3Hl+CBWjjN15tD16JspaPriY
RclRu5z/HVtqAFpTEO9zloG97C4U2UwRB/OrJniC/JEVRXeFZQrVhhQtrpJsRjXd4V4XZA+Kg6so
gOkifJA6TVVumd+W8yNEFR+VHgzf6MKIQuseubRlOIWFvRYmsB4muTHitEP5bBcaQRP7F5B4qZ1j
aqWTaIKnRBuNsOaCOr9fYBv14/VwoeWz4woTAY6NcAXoU1zrSRYUyRF968/x3c3RBED9Zpo22FmB
Dz6ZhlTDvpTMFF4hyUPoOZlAKVrsQV5pzd8ysf7WCzbPzoJ6kJGFIh4/HfX6Kctn6EBcP1Z9dfmL
iM/lYYgOPW0r+QeHOB5/hjLgGx0XcgbjilYZiB2MDhccD43INxjn2Bz9/YDVpRK6ks8RLdk7+/2B
ATxKZ9IXPFHEcGgGRZYPxe4N14mbV4fK50V1NScUq4Ci6gXPNYv0glfbUevIYFJ0MgVPNRK1vL/Y
feesqmqEv4eptKxMwz5QZegMrDVT1CuPN3UMydYxSnTamiLaeoXiokOy1mMXFZPtg/G9gpCFSWhQ
mMIonbn5vchdXfH1hZbS4grfrjQYcyayGuW1hu8dXCXXKNrki72SO91gsiczwZ9lRz+iWJD+LPNF
wxo6OqG7qDauXWCBB0QzgBXMLxzYT45Q8QyQOYDa6+scaIivb7M6O5W0gliOjIz13YSJd3Dpd0De
1T/28URmlcULUiVp3+qC93bfyqgqm7Dh1rJ+BvBWL1bqfDsq9tBqT15+1yP/6VHPWT3RVxRUrglW
FoVRIlTw/u7t5EcZ4b98rqLdA+YKqtnsprMSJ3Le5jtRyL6TiWJdLfp/8AKMGDw+S9xTBPqWOoON
2VNvahKhDQUycqdmMIjcTh+3BnVq/uXZLTuyehXMTcyvUsoFVqKB7UrcOtVPqj6rxie3FVUDlNL3
L5NEqB8Jkrm+86TnC0P0hEqIs8YrWl3e+6GRa6rak9DVvWM2hdRM7bqlOqnwPugr/gXcceoCcFms
52PZKHkrtPI7j1jAqNjKxhPE3inFTXWkqDPNgf54H7qf8VZqbek4+oxg33cFNkJSCw9elkNRLsFk
Pfs3lYcAVC+QZYyXe/zdMBTYqTQNgX2+NBAbZZ6IaYFUSfPV89yLs8d9zhalGdcWZgRsGqJEEZV0
h2BxDCddxHDhNWYXR272Y7du/BB070Wct4tOdKtAwFGnf7TCZ1i0TXRLRl1cRsRKhOu1HG2v0Ox2
Ah7UqTy8wpNgNwgbZZHFY92YHCfoRj5Un9XE7W0TFHBawqU1P1A7/0bz0tFXxkzAP6+/PMCBBaai
mkDpBQ6MMHBn4cuBMixcFWe2sozdfHDWSRl4SLpuQFmbRwr4PTeMod01/6ab9kMC69LCd23dqzHb
/GcowqjypHkwpPim6MD0s7UFFOFtxoxzfinIzpaDNN8OQ753+KNfTaVkhSFiEwhlfLeB8b0Ez9tB
8C2cghCwp1Wmrfiq8Bb3lDmV0egQMyRWYPwWUiTeb+b0X2vE7S9VhsAImNyBNiaua1O+Z2nZ64CU
EgYQG4GsppmO0NuIY268osytj4WvS6I2v1J5olPm+VXLpnzCuVj+U46ngqptdM46JDkEwJ52aGaB
NXak0NJOPjoqx3CpH0pDnjk6pCJVMJws2fWbpzngdUT2nOXuS07Orh1LxrMfSY8qPbavLDIyXs2s
tjYDH9TEL2Sg0QYR8CuX0HmkbJm7jkh5kEtwY6llVZF9lnYzmjAsTJHMxUb9q9E7TE86pbhTjyXR
Cii/E3lEv854ttS9jzOpsBMjYJ9UMn/mt8JiVMPWTUHBFF0MOntJ42m2AWJKLqd6KjaZEYqsdR7z
Afgu5cEDi5Ct1grdfAYhNAZIMgwt27BWFTHolKC92gd/g2Xj7udw3iCqMNQ7pJ9fAaeWUJpEpZep
yhK6PT4dNiOEddf2kWPy9qJlgqzzBqeUW2XZUxUhs/cguaX+fixT/QWMcDtEu88+g8dvissk9zWA
E6zj00/o29o5K3CZyqYuGmYCbaB7S4zIEKq70UdR+bBuYGiytXUNPAGJTJ5HcuVFYd1aXvWPy12W
4Oopdkbdy4J+NtUy7IouriN/JTRgorMvLdcapUYjRlvl860WrddG32vDt0LSYvCMy77GlqMuO1Fj
9J9ZzHfTNY13+vYnX28hO4TmsudPAnYg/s74nCmcjObZDB8O+3c1oG1xCe7b+pReFPJW6dfC1ZYT
MpfxzWBswvwXr7IYSo4v+DiOOBKO/4v7pYzmQPL0YeayUY+jz3mDlblqGchgMVFTtNtqL609X5AH
eekD3umhfzXGodV8vqlcxNqeyGvB2wE8kJnt4JncD0qgAzA00XIowTvAZfZwpBg2763e3lrF692h
Sj+HKU+Fz9RwAd4z3Tct78x6qC7JQf/jcvoVDuSAEfNHb84glZJpg05F5srzv+VPTomwINGqk6TB
A1C9WSg7gnF2ze/UgfXSFkfbZnVbLq9y5AO1YqvF7qJTPZlmqNEmoyCsZjBdhfMr3IVIS5npjv80
QDsgfsWSvEB5TFt8bnJcBRd6KJXvRTp/QhWDsCt+HufKNESgq0UPS9Mw63GoItB+5dL0P8AY8zW4
jdFaeFUHOjjC5b87cUJdU57uzNsB4iY3+QwOw/4NeZfYOtm1a8GmQqPFfra8naxTt0L8snmTPBVE
9//TQsqumtL2cRXj/Ckr4EcIRBwu2oatmGlRapnLk7VLc+ELmlkPxguf3Shp3IKbukGcKjnbZoWH
p2h64fdu1PbC1FgyuQ6jNuc0jbyIH62EPxsSozrY/2eA2Vtxl9RkPjDeShn+dtmzd8MRau2WVekd
spjORY33Foj+gEvhRBxaI/FPawDu0bf56t2UE09UXUHpIcJZVIoKiJZjdf5dcfLYnfllPuecQQKW
Yni59i2CNAHrTIwRyVIVudvH8kgoTbB3GcK83x2cgk8DOIF6pPqRU+bG36yhh42NFaRY5k6MsUgv
uBfg5DEaiUwhu4NkyM85CJaiSp9/1gBPzCTDiZfnBFDPwpxhkEi74/QBD9sMLefUMbUSqdH0RwXx
5vYLYEPCFxIquUHv2vrAclUNGsks3CF0114Wd+98XZPh1TAqmvIID3cbhI4T12JPRjav2QgMpk31
6wBRApRkPDk07budsxbHQbnXDb+YaoV7u6h21wmszDqsqktUolJm9ilAljlvdpbfB/NKU9xwoSsX
wVAkEuwe0455zYIrUFryA3uLI6ieGVAHscJMnlHY+xtydP6lwuDhEPtxCF0hjQHJgGoHAO1sVKwR
WEuNhtfE/0Ifsevnav62EbjGw0KbuMA0oB4NCrFFk4/QNRW8/qm3ZGnGNPFw24LoPhrZCrAct6vz
NjomQwOeFX6Ps9nPXIkZ9oDqFD/Wg9iDF1gMm7ncUU/0Gjqcq3pPjThNQm9tuZeEZug81w2e5TiY
dLWHqZc0cRIBKHFcWQCLjuHdRkI1OskAEmwocI8GjWcpi2LFS7/N0pmBEIXmGVmOWnbEoRxNNpHW
2REPXlZrooxJK74fpky6fiKwwGOzq+6w9OkDnMlAE178hqBg+nzt1V0WrqZ1PGhUn6IwhG8cNgO7
MbFhsKmmLxTJN6hom+Eu9QNMBDpTirsixG8TUutaud9dGFoKSzYGp1bPLq6rB0JYjq4R83hSdTxs
P0xLesM1F59WG3TpaQVnQu0k414zFOqQKTEb0x8dSGvR2rca58V3h6avpF8hM62SKv5CItNr/hg2
EXJHptShnuczUaV57D2jVP+s/RMFJgSUhDmhI65AdSBBYGv3j0eX6zoYvK0+VBGZhNEcm/T/KKpS
//Y/FtrDinAPFWkdwzGden8z9kppDc2+1AhPt/wKCSuYKKPXdDC0lMVrgeeSulX/A77Okl8zrOd3
3SPpH8RHFWzo4fBbZED94db5ObfzjrOx/UGOrZHvf1n0m3kLBMFYXcsO2TrVHp73pzoh4srL/p1O
Sbb3HqIdjMtLpRTfX1Q6AGLSWasoiT6R1Wdk0iP7F9zH86//QurcrAO/h/Srxk62wO92GEJ1q/8D
A4OiFwtVRmb5LR/K5bIComNJ3+01ysV3Vev/GjxKGdC0JPFLMH/9o/alkFBvnNHV2cdciBk3FdaK
EG2obfC50m/3V5DSow7kGGt4fiPQ4eXufgSxXdcu4cB0XNrkg0NAv5oMtg6QyxmTAfLxjXktzoQJ
tInLTAaU0buM8VH8b9eggrcFZEKIbhzXcVrXxApXHrkg8bN4DXCJUGGpsNJqkp5OkrJd/vP9cn0m
Tag1uZLGbmFr8SWwrK2tKzB5AKyCZD61rBzcuXRNts3ENS1FmXF20/ZSTkUS4WMafrjJZHcJIBAD
f29yEixaeVq1WsjykbP/GLaxI0Qo5l7uRQAoKHuh8s05UhrxkBm4YPm01/CRlCj52e0nDqVwpLBk
EpwlMUKbznR4PACWdQxX0fjy+0hVkjbFyqsifh7A4onr40vX7wgKs3L9DaDmXDqiSag6CBwPx84i
NVZns14ZEfCp/Bkvv9Cr6hI35vCNnImzH7jfTCZ/XZZ8aeQnbw3C6LINhSALYJUsnBJUMxPxiCr7
9bTtC7n9yfo4YMqXlY+2KmnEvtF/8k4zrSx7Iuy2BAnhu1NTzjFUXa/fjxOu4BhKynudX5seJvb8
i1nIZZdqXnjx27evaJQKd+iqH7yhAmJQDuBOwh4oJz9lPK0TKT+FGj8DoOPAfooXjmMNQP+dI5G4
Ja8GuT0zvQwYRZTUCxNZVKGGEIYY0mMCgUaORoRMdGvcF0dZadzBrKKYupUzTQiHyKaQs2cVAXsm
BwGyynS6p6b0JuHtLNNn/0yiEDyD4OCxZChdEiEyMrZRgABee/eCk6+SlukKdUjs8UZyUvIBQz2x
Rw6osLaYiXzu1q2hbwN8z6Jveb3NGjvLrkzATnSfSY3629y46S5E0X7MbtWGSdjZpKpgr2EQNAoB
0+4XVtKZWn9zl1UJ6IDN43CSMSUjcXAan639y0ocld8mqwrTaf91LQbYwzc3W5c+LhkfLUVE+Mkj
NKEZekbrHIfNsbEYV5NmB2EW9LiMaer/hRtK4y7/6yO31UZM4fFwe8HM5aOld0b/mxrLGvk7jojh
YtWvEcY2LwSEju1FiT94GBeHG1aagFFguIcMTH0mhovo+jQqxocvxCq0MBTt4EItp2PQWGNeGTRa
RZSS7YJWYQbg/3p6Ltg0G4UqKqrhJfTtPWdT4c5jMLDAtrpIr7fT3eD52aHlNeLWxHIUH8KRaMux
v8saLrl/ZaUFEi9m0arpZ4eVmmDPu+UH8so5TOt3VJht+8qz5qlE1q2T9RuQVHN8NIRtceXxT7mN
iFawkbUv/ywJl6zN9uwCwciJYIppnc6Et4q17jKRfRueZIrJjOvMxrFDhU539GMK0dPG2Q8CznfN
D18RvN/GtSy6/HoNCkHzvP8PU4oIHX1rs0eAFlMdzSFgs5/SANZOSBS25jkrLo05FANNRMCgp9IY
0WYNaZO4Yps3LgLvw0y17coYUYNDl5Gcqbk9SYYLBb5D0pKLjkx5ts8lAPaHy6NNint885VgiYoK
WYVtzlhfiTW+a4o3Bkr3NDa021cvE1StMHQqeGE7byk5gp9B2pGUlbj0PHLqJwVbWCMpUA6pIRQ2
z0xI+mY8YcKpg5/gm0gLRd5x3Dv6z6RNd8uOzB7Xw70Gx/ZmFi1XKlfnSr8SJIRCS8EQVIO5Hc4X
xOf+rfQVFjVcEF8sn5XW5OOBOiTdwC9s2bgd3xU6TXj349+0ySi8t+X4Y1MEbWeaYsoJP6L/X5Ng
jVdVNGC9jWZ+/UlOjdcf74/N2dEAS9v72u7HUHUehakim7V6TuYXpU8vgECVDONy8IYJEhP0deKa
1pPsTBe9TXDhMiDhy0MCLLHD7eLKTusDlOUI8p7IPyCSlCzVjmQnk+hy5kwIkkxCVREo4otyOU65
IDhzCWBkYmne5lSYlxSE3i4jj3G6YjUBQ1lUFdfiv888oVtISC0bCWiIW9wPZkNbTvKL8zFKqMLg
O/G0UEqEygiOnuH27dBNqfBp3NbYeeEQf+foW/sEMDGiZouRJu4HBxQygZjweWE+/0akiGj76nQR
zY6UAugAMH55FfR6J2LzTI2cwGmhlKQR36ILdXUsBMawnwypu7dXyvBjXVzbOEBBkvtOVE1W3Ter
GXuGtxKJma9Qr6zWJhEC0XjbDWAxqQbWeV+kKOsH7Ls8u0m2efwyXzE9+83eWj/wdRhigwt/7y7j
iPCkPjO2TDa36+Gp1HQ71ytCI3ktoiegdD6N6cthssdLD5RnrWeRddNe8gjq36mbrJGNfNgL+DjY
y2UrdzpJhe/btnT2OD5Ay0nFayxXVK9lIh0RW+ntenM+h6Rti7lSo4vobjp03bxIk8F+QHoBLaFU
GbzlCH4CU0eFu3RQknv5QfNIt9Mu1ZDqZFtaXu9qbc+y8q17DLopfdgahWfzIA/9gD+bdH7HTTMn
ypeB4NJmfmBZdSDBbZOnl2oHq1Ls8pLuV+iqWn6QdcRe1mXy24YXAN1REjgcaCDjosRP8CWDlxwJ
BwvARrNNW9T38LvIS5au3WURx4MLbTiAVTn1Q8sBrXYBrAWBEvkPHCdUMrD3nBY6jAzWOnSGTBSy
QR625BwyGzT8lxcMGIw/WG8IoG7CpNpWOPSMDA+jlooErAOE9khcu28rGyn/ELhlJdrwv1RzDQTP
oUl33fwoqMaJL73Rsd0J37FTliEmKwcbhDnlle0297zkQHo4Sie4lPHPl5F7h6AeK2E29s/7glsb
aCHdw2/JPwxDKdpkP9JqNhPJXgF9R/XXEl11i2bujSmpshSfiPNaI2k1b55ixKpf3hu3WySzqgyA
WOVLWHLl6AdNWu+8TeUo0paFaOc9gnyheThJhmPVCtYN9XLIikRePE09LMmTqR/7DgrVTMQ5/kBS
987YUoPS8vcotgU76ZCycde+bsVIY0J/sn5NtBXaLk7gWsnkfllutPDEXZKkQ317IuLL0ZXHXW1v
bsOVoCYH6AndhrTA1ug4LoyuyJVxDvAKc2x3KDRo+yogqJeu81XcAbp5ReaE4UGPFQXOmrD8Uzno
yKVHLeZmlCidW2VyXHQuT1xjjwEOgTDSU7dgqI83eGpHudL+Yc5BscgLL8vb4iOACh53zf2DCSx2
yzHQJqCoE/nUj928Zew+gQK3VL4Ly3ZGskn8BehRViEOMd81y/B06ku99LWL3DSxY61DchEfi5re
pnJADX6qGB/mQurktptRZuMxQqjN+sRP1v04kfTBnJ9REVb9d9dD0qZALCu2dkVQOkmWFGE0BlLJ
xEXCKJKhQUAyJhZCAVPXG1ssk5WH6XGWHulfjf+PRMArgT+vqx3RhJy8U7iGkLBaEBTJlefEhJOB
UpVm668Pyz3B5ZGTJpmkDdVKFzLWprIubO8lr949GsoBhdNo+vOXzvpYK7rue8Y5SaDHRshomzce
15RtbLgPL8Rt1J9deW8AX4617fdg/cZL74BxQ1BBi1SM40Fu0AvviKZXP8OwePvIH6Jj1hcdpSUr
bOPPE+FkzuG0Ow87qFmBoyEE+XVFrtynXXed2loZ3TdFIa3g/SQMsd3T1ZEjUIXLz7SiL0IHgQJ8
kVnrV3PKSLkv+3c0GDnnXF8E+sKo6HRlOXCvJNh6m7wg6mRzwPC7jWnPn32Ej7/SDMFYBoke713C
mypdeEk2/3K4uPfNIYhRvSp1UJ5MRI1vF4R6JZZfGfBGe2332B8UMB/yURcHezN/nJQzZz1jiChD
sO/AR/ClfPys6LTYOFJV+kF6+8kNPdBANgw+4cSovpMnF2i4EsfLfcxC3NtEomoHXIrGNod3lp2V
lxcUgyMR/CooGwue8UlTbojuSmMfmG8MSqsQFL2ojuBfPWJZpwm9wKD10gcl6aGlAf7ndMWnGpuo
Yhmq2+/sCxBEvmJ7na7pg9Xx2c8LsicahBMB4ppFb/693QvOShLj7Zn48TGZRUj6WHWzD4tVe0cz
oCJnqi57xkAkcRb7lZoNQ1ycFsNXIDMqpCS9456cdkk+OyNUFnLSOYhw2GuiMsRc+A0VpXLNSenM
ahI6W3PURudr+OWyhVr250IEvtoBJOoM/9AjxE6b37zZUbxZRyMlEEE7kzd0ko2xC0NF7Js6B9N0
rsXJtiv/+yuQHEJeF1QyJj+NMrPB0yjdrc9Xa0bzGfUrw3PtLdYwfT72/h5ZKCPmm0dT4ym5vnh4
na7l5AKBNoo7X4sZIeDUUVpL+V12nlvI9ryYwz418e/4yOpxsOS1kjGJCynsLhjSh58RenRU/hTV
CV+/mrcZ7jA4KEWWY8D896eIc+jOqlIMN3NYB0aw4DRNDnQf9bLrNmlj91eMsS0pKHjFyt4XzYjT
OvNMWupt+cpH7qhpp0q8oyf2f12L6/jZodVs/S/qWJwW3y5wuNqY37gZQPz0dWWNrauftdqsB+br
+plteiQ8F/y7mNC2tNrt58ueM2YLKUehZ4lJEjhceXeidnkKxY3lsyCrNP7V49D8UV1iQ8IMGm/f
r9wHZHZyA9JBfJVbW5a7gTUj6zK4gpQu9Bp7Jluk2t4oEy9sGpgPLkteei8lg/0gx2d3Lpyrsqki
8O7cOe1GXZMhfCeecfcEAGrSTIuidLd0yjoDPCGoRAjGqfmM4xMmck8Y1PE33nY9QpqSpZQOZEZd
8KvrAwmBTP3HOV4CjG0bbcHk0XdJWQAMl7lvEjfrchOKQqckngdBozH9bu13Gtuc296tReUv5IdS
o3RPtKIWFNo+mBeMLlb0tOJTqosC/5VJacjytfgqfj5cIiKL0OcODYWaDZf4ODmUJWKkI1uCbRXl
8FtyxZsm9rOIJFksB+i3rcQSR8l3K6Ty5RsdOp7OAQkPs6gI1wFKDOVvEpoXwzf06wFVIVOVax5a
U62X/a61i2Bw4WBVSig3tkmLjar5TRe4ThS2m5wFrrb/K31/5EXumEyv52R8uzbS2Aj6VFvztAVb
3/WB+qeiK39hyQlqoL7OPeKvBtNGBvJYaz5d7EVjDRCkF11nRURhKgwWpnZMCLeMh3PwUmb8ETax
+8OeRM98cZvHR+rkRxZEe2+R7zRhRfvAaDincyLIP7aln3J9yaUYiOrHVCvlpMmuaBZKpM3N6HLQ
2C+2y+hNS6XQrW/03vcLEqWd1WclXgvNiP8pPqbJoX/du8o6E+6lM50ipSiUjwXvVxRNUGICJ1FZ
fKIPA/91RMRQUIGXEAsiBPyUpCZ77MHXPHA/oNwno5TsUMiIXs8O8XsDldGsUexSKgxfrkM8KEZD
Fr0nk6agEQmVDWFdAFO3iFIidumJ3v7HTzdmdPTKfcfTEv7VXETo08fNrhACmSu6RFbtvuEjJaU2
66HqqKRZSbTIg4WVVkBa1HHEHoAxhg/dE/2FRm0IXHNPW0rJ7I5n+abDlgVBB/yKBbualSNY9z+U
eqarXRygovSjSeyesiLh0Pcxva5Te7ekKFh5hrtgHFi3h7v1n4SLJ/+NeJrq3IqU/B8AQeT4HmE0
9CfKbmaLVxTkKrtv1LVWa5adgDLLqkNh64HkrozZYf7GKlt3sqi8PKbnct86z0EVcTDoolqf2a08
hGS+Piief0YE420pM9olaYVA8djUwaIDifzx/ZM0HmmFjoE9XzF8igVXZfEFdJqDESST9q4fK/Td
C5oEgWbTSdn5GBPcdxszEsrUONGSlKnYlJQN8BW4zhztymc9XRYjw5etr83HLqnT9cR7ZyAQA4UZ
EK80z+H5zQSdAnnaMaSxDrL+ELcEm9AQyXY6KMaiDfhmfm7W7JeY9DErIRzJg6QHWOqkPyUqur6u
s+GKCrAn6hphR328xHerxg72PJh+5OAGzlHUpp/83AypiCNuKbfeqLdA1q/9LiHgYfWlIDcFHX6W
a9zomeR/7YyKxG7aJACDXowwMd3CK8phjcwg8jyb2kWurG71Wr8fFi7Hv3F9VPbJImDsAlbXu8ef
ejHx3l/64uLrCKPKl+8fGdqSNfaPjn5tOxB6S8CkxmtXX4lEbREWebMeD5Ec+0JNQjz0Oo8DCGnT
+yikgyIN/SHcKBRXkDcB2yvg52X+rDzahzzAF2n1FRjBEyOtajoIGn76rnS/GMQyOqVmWyDbsZMw
UvvcTOJ6jcfzFy+sBwAOb2j0Z7IYimnVjmwHSIxdK+EJGNZkhsGvO4U8UDtSCH7Tls8LvqEnBdmh
g40N7Cq2L4iCJYGEeyz+TckSfgjfRldKSua3OoVD07hTzhUOaO3fJhZpwDmPr7LD9UVbibQL2/jT
mgSXfU5lPE3jyPg8LBxXhqWtlakRQNqz6mDAaaCRYQVWqo7NHQfz4etOwZLvb2kd16ilRfq6mHQ8
6FPb6VfDrDEH/bSJtWaXfIoZ1ecCsTaY4SkOJ9/VwpI6YPJ8ak2H6ZVYcUL/2470uw0VKb0waa73
41qmobhPJG88wtRBDz+t5HzLj91zqkGoj92XHrR/wl4Sr5m/yfF5pKmcBP98cWt+ny2VMcoYn8rR
tFAS4dFvQ9P1rKODw2PgQW6oyHmMNhDnNRs280Ws9lu3qm5Q1V8D6VR1/8pL9bD/b5zwbFu8UprO
uZ1KBmKR+OgZvKqQYSXJi0akqCeNwCkh/g0WAJUISbqQU0rtj5/lij2+o9qCsxOvFrPv0kJQYcfn
/vbqmvcNArBmv/yoWRsm9UdteNyuGet+Ajjl1E2XB0aqaba5dJxSvueXB5u+lBILUeWST34VNmEK
8lJBHgD0p1UYmHFvIy9kJlMYlIt7BR2mT65cmuYkturR9k+toJMiBWpj2iaCBf9vYyG9gooH/P/1
9NHTrwGX/MgYiA4Zjw0zHG5O3wqzoFdbij89shhUx2mrFHV10VoE5stkY9eOgn0B9bW/MBXLni51
apd8cSImWrmCbOOo1K0AgxcQ01knBQ63scyyaJ7F5H3oKLOv6YqZTyQvEMKwPQMDx7Myz/Z14g7A
tI8FfLaFdUjG0Y1V1ATyLOmoq+8gW3m7PX7cj9G0LxWnXEsEG9TSG0fHJzDulg/vtO4v9vU2/F3G
tw++8lWs0+xqS2ybwJDwFro/IvI3UYxl5/QrTkh8tU/cnsZXwOZlpjM+WNsBQr9L2LoyCNOBQ/Ni
upR+WWpPZMJ+ORgBOhrpbA6kGmmY6S5m/2GcbIpijQcBh4RoA9RzS+/o3CmmfMpOwk3T8tnBIXXH
qwC2ottSkgpeUzr85J822YSxDqXl+5c6AdHW5/p4dE0ZwZLCPuLMQv/OcdHuwA3Z7D35vZHweJaG
JmbKMoigGt9UUoZdy69iZC3J7mYoXq2BcFk9/3vIyCK3R3iUMlFpV46juCyV0DogGsjoZyK7raPi
sABbXJkLArtrQyRySmqUI8WzXSfn99BY7tTGY7Kp4FFkXH3k6A/34IGPTEpWV4jF/rZpoIYIWUtg
1VkKUR4TFLOmzK362Eddor/+UeFdsTDodKqucrotkC7u/UVuPM1umViMf5/PW12G1Zz09b6Ze3/1
uUMNpUB5Fb0vzKChi+OuJMYi0lYbBVJWnJEEeZQfHyxsj24uincNFBA2RvMdPH8+QnptpUQl+O5m
qKTmWNGN6v3rrJl8F2XES1GERgdIMhJyyf+JJxf24GJq+teH3G5R1HfZ/UtuQ364NP9ZcDCYQPyW
ZNkFHSPS3+yS1qsfGA/lN1vfah8ubdYGSx4ZCorBYI13RXl6TvcIx0qJlXF0Zg2/5LtOruDw+U2u
uNRN/9OGdLjnPJdgwGPRQw70uyNzKfKm+TmIyjLShnH4e7DynH9lJg19nh8gBZuRt41d0Vrph015
aT5JwJYZo1zAaUr7E+hAjbO+kLlPy1EKNLyMMfbaH/LX9OG5IfRN297cjR6saPmUbf6SMQepL7iL
02tI2mvTlO+FPTHxvEt+kwceXpE/UKe2WHPxnHW+UaKem3j0rEsAiymKr62rfkWGji+gUYiwAQlo
b4t9cDCBxFr0cs0MbpgdhvhA51aGmHKqImjSd1VwJyW2Rx2HIZqS2VQcyrvGOfipcWYJJTPtF90i
UjYPqIHt6cT8kEWGqq0oLlXOUcEouOJ/ekNOZlWSftEdSJNqZVy07f2H53o5JgOuNHmwNzNXbK/L
INpTZZgmRVyyQWrufQqBbMEImdO5BF2OXFG7yJXkzUh651ETgEodPuU6+YirmIUxWDi46mClHzNI
lrK1oqAv6S+tmU8Pf+Hnd+vCkvEIDRRlUZ5wd0K9X5hujd4EZBSYJEHQTLWBQbXUSMmNDS7JIO73
1eO+RqJjIaYn4cv2B/9t/+t2z8Umo88kHfRTodiP3C4wtjvvPL0n0viV+K/P8XQ1nH/PyUlkIoKT
fXw/zS3Y9gtwiOFRG78XCnsGMyf3hfwtzx3DYZk9YEuKbBWLqar/pnDBw8ELOujoyUOb59eP/Gyb
SryUdbsLSJsXEGvaYyNFTpUDTeCni+8HAXPt9hELatkUF2+ERUZz+NBszVV867RngLV93poTJt6x
O8WnFVkHAG0ZLVKxx1SippQvIWLO4Z1CR4AgxSkTs9GyLB/0iDIpFOAchfXR5avEVbux/K+qzvKD
javGqUcr5KV7uNbPN9OwnZ44gkAXHtp2X+x410NIx/tab9nJD3IZ6XTSCrcNhUmbrda4a0KSN5ba
QlzdNJlzkwH0OKaepqxzZzxBVr7kloJmF9C/JB6iLWC+qPyZSl1tOrV3MyDj2ivHlheVqM1FJa8d
zt1WvT8jwSUH3OvxyWrEFcIBqs3Cl4o0Zm5kkrebXX+wLodZmJFf2GY5ydu31sjzghi09LDYPgfK
0kRSCLosHW7Ax5MwFieeeHI6BJ3Z5kihxtj7aYV9Bujd0DcVx/Ju6dr8Bh088852bhhHoK/uv8DA
orICgEYBnBSwBSD2BAE/zecOy8+K9mIBeO5eMnq1vIkkP8rcLWpIcwDTLJfFPU1266GKAbC1fVmO
xYV9VxXDgH6Cdoz1uQOAFG1MGDM7GbVeaQJv2bg2WjYLFyMdcspskD9IsEXaIsPSnpb3Cg0jOaS9
iqQEPA5UXwN2ht8LM33ETZcqLQ+uRe8SOH+are5ZXLC2B35KYB75yNqstEAsRtp3eIH63TpHMZ/+
Ih5gWnoyMur71PfSD+L49XBMHYWjJDY2tmfvJXg/Ex44rAPMkPgtsHo8v6re/+EoRPgThpkqLS/L
+hIjLEX6N351k/ovKVbSoNxURDuku50nTfqdHxKXrpQ36QeaU2yrG49U1ITNj7xHdwHVztOpd1Z7
Jn6uku/9ISIjvmzYKi2KddEYHGuA7ze5EbCdnscgYhLX9FT8B7XNdZOirqLlRJMeRFuJQAfoUSST
YhX1qh/C81wlz+9Oxi2xi/FeglOrzkNO7Im2SsazQ+cn8F7PDqBrYiuBYbwDYg2Go5LMqCKkvCh/
KtJxH9r1+pK2g84bq7NaaxO7RVjqq1oAcYZPc2peXmH2ec6rv7Xu5NxlhAlCJVqo+mjCRgg5RoQz
l2VssaFLjzrUgy+IUWxn7vJVRswXJqEUogX3+pXu9a+QFPNzmniaqDofKXbVg7pBtxTE1g5CZU5x
k9oiJq80SAlL56OM23T5FAHySzg3c+mLF/E0nL2/nwxYs0u/vD6GjG91ddnCl0oP/TDu2jIa5fuY
aPIXxG2RVh9Zm+LZ1BR8vs99083CnHntKmWM0JcsQk4fSYLoxeCRnyqnNYGgYP5/WncXV1u7e5WL
swzf6mXNxB7/yncrLSAz8niUGUXFAWh5mSL30sGbLTfML4Hrj5WDHMkyZumT5gxbN9RXGUeNqXKd
y0kXuG2evDppVR1MF+gX2Ji3L6BL8qRhjEh0Rrm10GGQhusKKhx1vzzFnQxLGLPEgqz8RU+JYopK
Up7pUhwIrVvt5JfkEmGVS5nsUmFor1c00Ke7MhMyS3/siag+lg82rerwAWvvN8WoBpJY4hYyGbY5
Yr0yUnAq1d3xJLtwlwChnHWXafHUOBwr+4numZmw405S7S28ozGrXJhoYd5nIKNXWMKS1UTLlN2L
HuWp/V/VTxl+P66np7fhDIwu/au+Odhl1cooNMuWzSwf2Y0cf5x8GxTdWGpzhPMsGQDEXEYzigrp
GKzpQsI2kkP5E7xOyfne/U47sO/IcLVlLAqOmkaqlqwj8BKBr6Xwh4eakYL3cPv0Ap3NkNFnEkwt
c7lD/CH1hQLZiMxpy3h+IMR1FtJ65sL7zxxXeSnZuKIg2uFn8Zt8lEIHPWUAji7Afuwjc41y6M9A
HaF0KGj6hYhp1r1G+viPDq1TZhuE65aMKx8yM7bsAgMhvzM0J9OLGyAMAphMCaDzUqFwSHymRh7c
byGFO2APzSG1D1ZEp6AmqzB2LinmApDSxX+b/5bYIIHr8YHWlzcb/oA0vJ970LePVD/XuRTnrtYO
QHJWyZBP9k8JUYZxqQj/KsowrCUEoYDOzmrGGwNd4FO1vfVLTR+nf+onTH15ikkigZoxNDrEaujE
CjOuAktaQqRoItFasDVR0jjgwd2l54n79XYfn/yhGR5lUjcY9MTXAKY2J1T4tX0UpdjccQNdbLFH
5fCNjRePVTzVe5FHSNML1cLP1zjqUUeR/DsNba9t64k9k/wFoHFxYRph56GNNewwu4VC5DdzI5Ap
ShgVZVtlnhJy4i/uY23pRm4esem4Ehs+zdufNGirqWf9fWsIPd6AwU/8CM41rkFPC2w2anABKzw7
92iDRJuKbeaeEFXdb8Bwcdk8vpzNZm44VbJfUyAuLSE4x9vKxYWKfQV35j1sTYJkd2dQRpX3O2QN
Kjc2I0H5IH9eMF37WfmBftwcL60nidZxaWUbFQaGJJV5LB5WUkxYn6UlhHC3V4WfqaKKKxz3W73k
ePCKl7QIS161BYlovwwC5k2MvXiCVkHVaJ2aL5vGVAVWMBWKAMfiW1nfhCRNj7lmcxtW2YuNHgMs
I6F1+IW309vwq5eBxudBe5I/8szYiwmaQzMPoLuuAx/+7UVVxEMn4n2iw7b/OHQ5F6ONjSGUzzjH
qLtSaxPxpr7io/aDjbNy6zZs9NFqiD5nZvYDpuR6/tvTqN0SwH+cOpWQZ/lHy3njendm1qi2q+/7
kNfLzKf0kOFsI2v7JHiS0Zie2KBYNt9RsIaqHnbQveg6ZNyizWFbaAWgpZAzb0eM9VGUqezKgd+A
Sm/RVcfTuiwTSepqL1nNeDdGyxip1lqX/ayIjC5iCguG5CHm+DbKuD6gy+er36BAkjTpHbXh7Iax
eFPq30eMPyUvN5t+P6iqrUPDhuYjX8n6qTDlE4mX30PkI9aqlmzTTqShsmU1YFRtOGBur39Lxmn4
K2EWn97YlF3BgwuhNYgUBiAiaJ3MLueQF6GDvfyaOXpRg6E0tyNkP4xqL3BkIcjTkOUtPFINGkzy
ZFonR5tQrG7rWFVWYfQevyBIF9VXDoQJ24DLlUQbuM3a0Mn2BakWxjVo7jLkRNJ+9ID7v0sUzMJv
7ODljw+HHwybRB2ewo3xiJpjQrUfIYrkLNiY5LWYnS07JZMyXBEAiuIWFg7/ZAvX1t9wsrGUB2Bg
GGehyXaRejFLZpR3IXsV75XFJaY4saHIxLauviLmCSfRLFQmIfxVzq/CxNkt+Sdus0UGY9WJne6J
WeedApofWtY7mpn2rxHJGqOcce0LGqyeAU2jJTGUEd8VZ68lEWNg7IWvSCc+moZEINSm5cuPIdlf
t7hihbAl8txLdIRDNoOMbMgfkVrC07bzTrXw9u7VnQEbyHPBD8Z09ihO+C+nD5SMPJRKWReUzSql
RstrvoWaM2EsMo+bV+d7r0fChgJfs2T3M57GTwqPsNIBgQzhBEV52P7DAI66BVEGx3cSYwyqYlBO
gZZyNtdfDD2F3+pBdrkP/fmiEC4gYjsG8qs5R4/tjIKMyYiO4XcMNvJ8LQ6DFU6Sj6uRRgYVYv4L
6HeqV63XcG0SNX9TAwbyNmZvnrndSS5JVGiaHDKunxdSkdgyFcNKlZ77230KvfeWIO3Tyj3mo7GZ
zVP3mgmwI6f+zLVMvN8j0/e6V+TZlrgpXY1r5vN+77gZGmEYvt3VrY5z8AzGjlwaXdzBXvwo+AMV
wkFviYKkf3ml7YWz93QgSbzYWkQSpD68mKXTosLNzveMOLZGmfmhAFD6dtk+HEcP1xeu7+P8X5Ug
zncbS1uQ7CdEuMSCFYvVoSlUAuO/06EGIhS8j4vil+lM2s3ZhBKxmBkPeXlf40vVe6MUp28iY7SP
foSGh+7imsP/xpoEkf0wUHYLk1kC+/rnMwbJFHk7bCGRZEGWMo/CMhvrZco/UrZOR7VD20HT1xGQ
2U4QrB0ivCxSOxbG6SLKHDM/pAYYw7PJ/+s79DVVCMHlM0+LK5tdWoEaKnONgGo7lU6vuzUtdZyf
euHieEkwFDudFZ7616gWSM5EtrJu/ISughCGAHWJWx1Kvw4A50XNBAGZ6OfCHH2+zqzJEO2mgaVu
WGblwpenzyIMm8arfpaY2IicRO9Pm9SGFfce/gJuCewq8MJWqTvhJa36csUAPUuKbJ/JBldmB2N0
lWD6AVV2C75uNfzoB0ONS21kHnKivlJgMtt1GIpgc3cF8kwWrqSyF01zuey3CiuWTxJQKDEKJAw4
NcR3gp9gOEu37gNz7hH1bswwAzCtOON5DEf969v+3dqHmHdL12Oquuodk7oH+cbjG7To6MqGbp9c
QequaMyEbPMfU+/yNa0p96Mf5d/G4bxQzZVMmbyx77Bw5V2XAyilwBjH1rQed1CS1Wjin29dOvCC
tgMkAJzUlTba9yVhopGUC22GqBRKDUBjY1rWHaiINzdttr32Z87MRyy6Ji7cMRKbVWIDd1nYv09y
BerMgE8R7MYEBcRr2ZTkhlW0YWG+pGVUaZM5Z9Olx99CKLpIcx0lG6ZCQZ0kEV62eqgWuV9aaHSF
+qErV41J5+8r/spHKBrDCk5iQU5+BR/EAZrCkBwfTMN9qQclNOmaNrpgWZ6lJ+3Jx+nESkL3Usc8
F/D9he1HZKrbDPEPnbrln7gVzMevZ7+mVDnVOCqKV6f/wv4R+622HrelSyoXdrYxU1qoWN53Am1G
GN1/xtsevhfscjTGlolDdaJn0XuzaCZovxrqpuSCyGK1pQ4PRtwLXvdkMEJMthjlkn+kTW8SFiW0
QxFYSBuKtuH7tIqCP4GuVSw3bXAPtZ9jWR/ijEHS4SnoDtRrXX1fCCLgVHJZ/dJ6IXZyXl8J45VJ
GsKILVGolCQuu94rOcaOCmWpGOgJgRCm8jo11nAKOsfV0rvSAPhkNfiKkH3veR+UkjdliKbGI7hY
+2g85zDYy/L5fb20GV/Fo3ugSv93vTESBt7HiX7vMEOp6GkEQLYvcIA68QWH7/PHBopABrVob0ni
CWdhwJ5A55klFU6THZt8j1V8pv2ttcvqz3LSmdBJaTjUN893YJDTRKoVQiV2NYplxWzicsQFif7T
RpS95b0a+jrRpcZEdSUS9gGl+rhE/5JwY6rDDNz7yMCA38ZiCuw3FPayfhcJhHP73NW0bjRzLcyh
sRN4lyFkaMckgKwFcDKUX7jRbSInqMLPYxLPKCQ//3qgdqbZ+VzNa/S5ug0p2iOc2xjgq5QZgUKP
K1dYt+QEl3xSzeARU0ynbPiEf726RQhicMdmemdRVLNvmMxYxbWbdKKkgbCd9RJ3sbRWQBtCoOdt
v51LuzfjZGJdTr9L+uGyntcEdM2gKt2zoe/UWgxqsOjPPWwjAtnoV/02iT33ItxSYlqmHrGWs+Ya
MdcPYmTJqm9co+vyGGplJMs1RPjXdR9Aa5K3Z6rvL04uuYy/ULh9y2u+IpQAhPZqKOOkdHulkK+z
EBzIEmR6h3bivhqKyD/RQLUZbSM8zbIgcLucc4zJasgxPwFtnMk3+X57D79OfU2Xp9NKa7bCnM3C
teO3A6D0k16a7oztRsAie0OJPlsZ5CyM5g867SdxB+CQFqhSV7i4CimnO/1FkaDItbN9hEcuGSif
SYZkIZaZ2tvDuVzqm6cH3V9XzrgevDhWkUwYGgCOyvyOP5TWnF9dtJ4FhTXquUR8Cy7CjVM5u8aS
baM2opFKkhFixP3AsroIjm6FwOA1o+1QvNsijy0RqDbDglrbxZwzdVeiYCrpm0pu9RTJvMiII4rj
JcdefewatWEiljedOqy1uDDpj4XGSUSTuwMb9MzdEsQSj2JzVaDNtfUT2SUwUR2kP2DNI3pZyyg5
qQVDAVHp6Hf4204ftHjTAn98mw4za5hWBJPJhwlFdy2cB90JFJAmx8tPz/Ka9hXW3O4POhhVFDi4
55ghCa8NoxV7mLt39GjPEOKnAUW19EZHd99j7Eh1/ks6PCKHAyi6fJY9rCsfVBMTCJwwtwKcKuCW
vxTX1Z2T9nEVhbq69gE1p1RC6V/leX16S7DLNmSW14GzBcXYC8/OJlHRDsuHUwaX9xErusLsmQ0D
cbBn75m8csUldYLmhPlEsMCiaw16Ai24kPavalBc8qytjYDH1qgXQiIrN9NA9x4EqRhMiMbytG7B
nn/QjPBCEIofniTr0kvTan82qmb0+IQHXvIM9cNHlb3QMym9HLThMvTsEyFXxwfnSWJCZzi0rhkJ
c8CVGZGDwVaJvmdCHnl/wQL8vL8L/+vrurWWSXZNAmxkHT12p7Z6YdBfWDWyHE69pJshw4OTfO48
Au2iEPqDTlFAIsXsdI7mW5ps3FavD3ewRPWN0+vTwadFbeEuBvZfGEnrum6Y58gqnRjbLuSFZAve
gEwtWW6A14u0ZUVIZkeqOrzYPMsQY4VZ5zIo93Vk4v8NjciNoK8CB8UQ1dfOhXbiijUYyjlgOMDu
8i94YCUnPOllm4oqmsb90aj7YLTYPrBecY/j2idrtZzF7dbd0doAGqiXxJ8UFeiJvDQjzNT8r66s
gOC73Pc+194JTs+17a7NDUY2bp1EJ+vqBCSYB+nlPjM4zAPYYKwHHwzVB5b8fn7ixji7FktI3dOc
hFReH+DlfNCITK6/dgKFFlpNEvk5yJdkhJA4tweUlzu77Byld3qq2zI300m3AJXfZPMj21HmSa4t
ipxS4HcxF6YdbD/vxjTm9AR08obnby4JqzobnxyHBA2JDMz93HNVpA5EBbOrla+DvaSyG9gJheg1
7au5Gop/ixIyQMsHs+vUV46YJm3nZter70TKGKZ2XRBNFANlHkcC0hGiEDvqPIStFA2YR5vdCn0P
tT4miN8OQnpQs6Avv4mtVMfyVj6aftlG3SHHc/raIbqVLs9oj/e5HdnwLqRuyzjqX2IQHjIv8I3l
i7CPgPNxYSV1RgOPgLZw3iaIxt2X4zcIIgudFxKUegwfxClPmivfxqmXcbAgiqxFiF5PdvfAKoyq
mUtww/2TltHVsrtzDA9UTW0V6/7OXZqvOSlgaODkpPFLnaDAWzaNvuhW/9d5F+oSamV/s/yyOzDH
RQnx4R54DVefKDyx37j5/xaR1dENM3MD4dAUu4e1B5V6lALQyaMc2acOIvft4AXXFHa7WuIAqeAz
R1j6yJSUu3Rn+hc00LvBF1ZxhtaWpwBg4fgB/C6sIhGCW6aR96hwFFfq5MHVR6KmPK228rgTeXU1
4fQMf4I4RhAWpGq4LN+R2KXkaBo1uhBO14NKylIMVYlWpYz1e4oSZCpUQKjzeQsXv3TaluuZVryQ
XccDIeX4ctMR6DvkpdzGPkjyorvX+g8Q8kr7OLgzWt3aLK4u3jC+FGl8AOI6JBDUVoIBpG8mnJMf
dUmyNlU8eCv9CNAc7Fp+1bb0h18qO0HR6abmOJAXsyvl33LU8mimdT9Fxr8BYi3SZPDWaImKZ9AD
Rdv2fDpNArWxFc0Rtm/ReH6NrMa12WFuFKJLY/X9iufspFd+XkbLFFZi7bdWNuUmG5tRxWgCIdyb
O+3cmxjXgrUbJPAkWZmSMNVo42yfwwQRfs2cqMhkmzXlKL5OOJzFLI6Zixvy5jcRQOmfF9cnh/oI
6nH0QWLHcaHwJtQiS9h1jp83/FM4h9Y5ZsO7IsrNV4vHsfH4sBUFIwgRpIXERmcxk+NyrteF6z8d
nQDT6b0nzpfehSKdixdPJvbESnQclS59vdvOL7QL0A9Bk+Z8Z48akFOsJZ/L2jRt7R3yct5eecm+
rW/MgRdYHF3y0ccHxOPSebOxFhQIN5T/FgbFNaaCe2BjAEcO/fu1r43EREt8x9ktV5ixE6To7on/
MV6OvymM4CDgcabl3/7RK3UUlKyxcweagIYv/NB/XsxxKFIRuYdJT9cg2do7aYIpe6El6+9B3bMl
it/LlmFsSBGPzjqyzfyBmnCrWMvdgJ2ESaXvAl9c+beL7PPdhXpVoRtKfc+sVQbNo5bQymlrRCfa
YP1sjuQvBKzHtQofwMdcn18Hl3ucsXAWreQpauSZLZJ38/ylFMZWJLqg2O1gvCbn+nDUBtgh5ued
Ky9DTSfOYvNNQ0ZMlkq34di3rlewDAfKMjorkCGW7Y973UHd8waI4ttjTn+myq7PLxQfCOFF1WLk
dLTfTpT0xCEFovsiAcTsGdCLl0l4jYZJUN609vGmp30kFpoDVXJLqvmosiWqed8VDolr1qwdFX0B
xCKRlsPtMnMRM975t42Dj14uB5EWfbB4coTteepvJc4ym7N23Ua4lcm2GMo187UavG2i46iYVORI
OcyJpLVbcaRQby6Vipkq+0VPlG9gt6PKK4PQVcr/sp6YGsWuzaGUsll9jcOYYQ9OFuNg2MjARAgG
F2aOZ/1xbxOSCWpEPLKq2DtH5v4rO5wTw32oaXD7xDD2OpGEED87bWR+/ZVoPFcVTJkUm68US5oh
BtHREltn10NUDJbQ/2ceJZ3glsFutcF4GVyQW+J9nz0fU389g+dU2oDZ0mAhtjEWj3VofSMI53Fy
lD2QOysV95xBPpdFzHFBa6R1gJxjrOHH5ZYNWFzx1AjssGyqmX675IC+ohR/PeBMgouIR4raGAgA
aGFmMBiyTJ3NiZ53Lkpk1yN4Clwvu80TzJw0QuT41IKkyH5tU3SNtKh+c5+t0/vpmE5LBZ0ESpG5
bTCQZu2vZBvmullRq8cRvWrlbMGCSQP17zUh65S7DV5r2eYZIwIgdgooRwomWPvp+XJm9Da22V97
OB2HDduQrvv9AcIN7TRoNnQ46hakun7iC6sWVfhFIoS5rew0x+T9lff1XNuj4c7LH7gQxIzCBSp/
8Z28WMY8UvJmI1nKoXfyCfAGBInNk1bGjSUxI+Pb1LlRUvYj+e/0ELNu54xTKBvI2eYXSGGH15uM
/AAPbDdMU1q8UD0ZAIOATlJSDClIv2iZNk4uJ0x31HNhQEPpkkzD5mKXylZl6a39Rtq51MY2/S25
w2FhiqoHtxliVnjJC2A6r2fNLCOQ4djip492gGqBkdhfD1QWkE0zhSqgz7Mz9NJyxW1dkIYKHDfq
mzleEiLM7LdhZn649/rQ9zXSxns9K4IKbIknaXYPYcnRF6pTdLLv2oO9txxjRd7rH2ixSsJAfF0y
PV/UKi3HncHLu7losEkYvbeLROFCzfzsvcO7prgxcsMf3A1ummgNIw5Y91W5WsNXdlV8wst4JNzl
ezL+iLjHeYBm48CHnH6vEkiNPvlUGHNnVvmb+OSs7ZBToPuKKqd/fSHK2QAk6Bo+vHuW54mGCNzx
fUXqX4j989JP4hu4zTKahLohM/pM5xTBkuM3da7LGPdkeQwYIXtOOYUlN+8aZzj5FibK9TIzie97
LMJSdGKBVkYy7O+dMrWn3tv0/yR74ooPdJACvIGyixHNDU56di5MlVy2xp62uWdhRB9T11YN6n6L
lJgWCOkwLZvINm9yjjlfXp4YvhCozv9Z6ndQO4/h0yP4CqrqyYmGtYE8GoTK6X7hdSdDt+yg9jo3
9HNYB+SBAYRFEv6MqHvaY8EJCytl4s+khTRJHKPE1z9/o2ogeS2RCFJXkQTSNnCu6O2ltc5A8XX4
IpR5WbgJPqSxBf486uodXd+6IhcExgrLLgTlCu+FxPWQtHfkx/kjzG9wX9vJmZW0T9JpBoDKRpNf
uHZIFD371N/6aVInVAKgroyiGfu9+hqKzIVuulGSc8Vdlep255LqDO9Xl7uH3Ztj5jqkZbeEyQwV
P7zpsDYRYYGtFPvani4fDxmB+w1h5jprjO8K3SDTcRvOnmnL3RGL5PhHQNg6w2KEOYnko+hKHk+O
KFGv32O18hbCnZOnsDAmZhbVYt/7zigPnIVmzKkF6LMyMBEtQup3GjoNw/SBC3kAKnu31gdk4//J
iRMHn5pHbwlmo8TA0agJiAa6CRXYDe4uckBVMsWlUVuZkV4jvrSse10HuZnIyDNW8kvVP5a87rLp
yLIINWj1DoIawh01Ccy3lRVdLaJIDZiRfx5+JzzDNkxb91JMpTy+tzKYdRtD6T7GceQZThwBORoN
puR7zGENvkkmUM+aHbEPB+/1GryFcW0O7nI0cftiQsakNfGHSZOiBAOTzSsohDCGQeYD0ICvvluR
5l1Q3O/+M808fybptPlify/m/rejy99oNM+9lucoSqvfUXgrgFM8nZQaDIYBD4L+hupuE8gkaktL
T9YGnKxKUcYPhSAB/v41E1zD80/3N4zz88yURctIX1bKU3tvDvJ57VowHXgcZHTj3xBTtYqkocH4
Rp4QnZyU3pYesAUGk5vVMqkJogVIbRb+nbnzNNZD9ZASrYzUfh03LJunQw8po0A+tK52nCC3od83
rBEsHaOJbAb2ahC9IIk6v883Yj20UrrUEwHPVMNl0W11C6t4BHN/jAeYpVSfD1Q7rf7YYGpALVba
ve4aTfiQTeaJYno3BaUZf1D7dqPzHOV3fKHOeHvHCtMG/cwo6VAVVTmuc4yu3G74R4OvHt0Qhvxt
akTAqGOxaqTwuLNXghPCjnhwi7qUZnQJK71tKb4m1wITtV0Q6opC+UG/kKnmsE0tUxbvKnOkM4cH
B2anDJiD86rHm9SvMV95F9hH4gbroXMzoZfoC7DQsTJdKjAADMvKSXdkXmJe7mNKJ3NBnnybM1ao
GB0H9AExnvBI0f0QxjvctKkFQGkP+S1L9Td13RLNreoO0W0D8m+cm+Ood8gBYpmvU28UhSPeEvEr
RQVoCMXukG3KLs/3j5DSrmnVv+rQ+0nWIAumSQxo1Z4wW3Rnx47JOxq4zC3D7ZYez/iczFSyADcH
t7VRPlz4XGEqzWVrwnYdA8MrmNrhIrE2bVNCUPRPlc9oXlNMrIhp8tYP76dBi4aBy+bbKV3jpQCm
z6Tv2xc8bly9qm2xLfhYmu6+ZAzVfDGunqMz//KPDMc3qOH64BPzfTeclgXE6S8bUPjET+UdFXJJ
98EH2VXkcgNim7Ajhpfu2mOkNPzvNvo4WxAsY34OLenW41KyZtmL+TnlqaZgOhupzBsT/+IKn82T
wSaWFxDGATywIvLkpPlDZcQhpTfr5diFskBgPBqQbXbvR94sP8e/NkYiRIJSSRs53HpwaGaeAlTW
MuQP9fFsfkl2SoFwr8XEt8sku0Vf6q78znqaLO5OiKrXSYDrUKRBG8WOzLN2Q2QBA8NAbl7cjtv4
jlJml8Tl5IgTk3XAAV8YwJVMEvC8O9axF3G9BRbgmFx1P4JaORzZrYd1uuJGONIiFRW4xh+YAECq
p5tPJfU7ObTEYlXZGezKoOobn+mBq8FOV0n3IVLx4rj5YC8hqi1p7MV1uSuubbpCytl5dvnME3Bj
CQN+b+528IU99fXT70tfm8WTdovn93x7eoDIMQ2Hd1o/BG7koAtsTq2Nzck885HKcIc4A25TTqdb
MJ//NsKujpSuP811TCGDnwjcb91H0xWwZpYzLqiUeYmQaTPu5etrHDlwukFWbWaA91HBNxNqyZ59
3rwCUNVWwPs/TfMP5uKBuEYkmKaCi7wnZe/Am+CKiNYAs+JnyfMlca/+r6dkPl4VmYtZoM4LIo1m
AkgXdAbVIFI4i611m4QV4rPGDC3m4lzEejScPvi5RRQyYAubJTNfIM3FawfzxKt+0E5jAp548lme
dg12EJ4HRXMamC6OHzvAfNBzJqmmh1D/82C8GhPSWOl/QMNYLAqd9QDbPUbOOQc0U5uIIHiG8ex1
P8TREd60xvrhPdcnRVXPFU15XIxIJPea37WEgz1HmAema2+DcYIbACN2T+7ThCdzu+Ht/FJWZtbz
PiZs5t2Tkx2TrHrvGtdVULu+1RzVzDbWNuJ/RAMNKpCNDzYtgjc52yrSuliZifd+za2O8ejxqksk
0ey+WfvHtj0VQZc/aT2t3OwxW+eN/Hs+kzpxHZo60xaJWNFy8yABcuUuLBjFMP4WlKIZK+iv8z8j
6xurbGPYgeO6khqZaW6/f8lGNqJB5AJGSPf41kXQ7C7QCfwGfL0C/XrNrdVQFjzomTl4t+k4j2q9
BJrraORgeJhCjGZsUrJgBJrzgeXkf+QpvBsH5keF56RNQ/I1AuppJHUf06Qqft3T5tgJsz7SIjR4
kF4ECyNVijTWiaqMAHyeTdNQBM2fixGZWaeLhbz7RBkObqeLsK4VqQwa7ojDvxHjOsW1UrjbxAxM
8+lU9Yvah29c+7/w6NFFV5OR0bC50pOa9tHhvvIiRfVLZXBNePGBppCORi17/mActuD41skSIpWU
bsF4RDvYuxlKWkdKm4PZSaJUwPd+WFi+aKk/mTxqZJwRwFsiUXZiMtxOeS4cgvN5LQi7fk+t8a3B
ySzPz1gr6nLueoZwo01oYFwDmbL4I+wYSVOyyiibTr5Pr/cNxZ67OMQKZ6XHwqJ05DY4tHNmgwR9
C6ACZLN88yYbmwIaPRk3anPrE8xd5494b5T7nk9guinkkAvVZ0YrYv2BZIttRyRrStVttIDLLwtq
37cIJ9TDUr/R6sO3oSRqcdel+QVZwzPD10uCjwAjBLpSO4kTHD1PulmglzzK2rxGjOgFlP9R7ikd
KmYc0wed+Ydo0SiH97RFT8fq6+cLrOZroxvN72bTKJk2EpM+yTiYWvwbETD7RaG0iGAhwFCnDv4b
ESamcmlkGsZRaJ6TtoDGFyBmXIGVmT8IfUPt0KUD6D/7p6hwPrxqfxyU+uyfvzt1+p4CA0jWRDTy
sSmY7XS+LreVtS3shvBueodFWNg+kO7kPOuyZLkviT/WTdrVxXIWuGOANJPzsjhZschp4rzv0xCr
Z5rqg2WXboQzkfZJx7L0ugClr+TfyiMvBXjuxAKzIuPXGWu1kmmzj3sG9quSkrl40Ofv42mTxbn+
AHl1skuFquG3MjL1I0UK2XdiQS37DGG0u9HkeoJdivoVgvTok8zvL7e1WUDR92MbhzWtlEdsXB/v
RhY8l4bzRDPbKcWkMDFlOeo/9fTxM8fMz/FR3/FsyKPCOEGY+TMWsF3wpn6TVmaMoLSrQJfZAXXY
GpdqiSwcHaj1JJgplOsIWxTG9qadoSkrz1q2jD9wEiW83O/X2LiRY08IjbpgYIsYlcVlaGcegjr3
lE9sQOOXY2kY+ZLWYjIrMud3iAYnf40srZGu3I+60lGh0oi/F9nIMYsws6nx80e0xLZLIoog4EXx
fy1JcRisF7eS+daM2X6E2/pULSjDstiXEPWlTnCClP8TnmyoWzR9aL1r42dA3YjdxY6KPDLy50r6
y/pYNvCT20xvUniNjXJZzgJRKXDjRIN3d5EZdFWWZxUvVefwztVHXUynKJ6r4MLimqfB0oxnxpxO
GTeJp3/akEB+SC5TusskK7j8hNAyo2pAic3poHX1onfTbe7lG+YzlrvTg0KP8SQ7RuYP8Wfh8dHs
m90rne/5chGQSRHRxzZmFP6PhYQ6C7quDG0HOLfs+7u9CWn7m9mmFJwK0YVe/TdF17hWLaitgdtg
z+27TDgs3E3TGvwzWK99JLxG1DSjZMqnOEA59AGUes/Liu0LcLHbxPLI0Ij+RLjb/0gYs3c8c1HF
dyUs/Ad8OlHm9H1KMdT1CVRv7sTxTvBdpvM26eifoiAn66T34avsyYb7zJkj84cJhIT2SQ0bqwP+
RHPqNa9Yvr2VmibTm3RBpmITvRlAb+zdRR6hlnvyOWxKX9q+wILKla7CAfDclx5lOpmnH8YapmNl
UTqFg/Z9tg80b0Z7ARlTwg7tr4J7GlaWAihTmqKN9GmYQCgO6rzmw3HJlt5lUf+VSV428OUUwApF
4PoDUCvhVUCsL7ZVHSOuH8jn1xJ7b4TM0rF0dHhM4rEQ3z5qFbqd8zZK/Jv+ZkSuvnLDskNl7tgC
zHOHIUScDfdc1G/tEcHzHQC9HqCDcm04uuNG7hqzwKqwmS4lGbhSrKKoCb+oA9vjuiIbFQtd7Xpu
dHe3VNcQuyERk+O45U5kUyJluoiadIBVR7+v9Ie+KZxwErig0gBYW4G0dc7q+XhCv6U7McHw09GY
xOpKwpt8nOn2Sc/A9QLuXxw2W/2UvX964GRJ82X6ywZnTDlKDw9jwzSQu1OMji2J/VapAfknie0I
Zu3lmts1rAJSxhB/2JbeQSNkQRPVanolXC5//R6YVToWAwRrqdzDjUQnXWYzIq3WeDNRZX9vcAQ1
gQgpg/AUPi6HgIOsZy8Vu1X3X4ZW3PEL9qsYyGsX0Vlu6FMSHTZq6gRf4am0Z3Rhjg351dR76HKM
D/7wkxCH90H1XBtCeAHBAN1TYGfwQ5GRgAmakF+RKLdS6jRejkddJY+2vv2rW77MKmUQ/CK5ofKP
EB8W+MHh6afWEfO4ErAgHqUwLXPKwcAM2y9h9xGHUKqX5XnDEro6NbTJYaSxQVNs6r7fKo3YWYzE
Z18+B3V7fP7hfxK0mlSDYTCSEcbKTyPuEAkaqwIxSHe1qAikSwPEtE1hDKp6qYRzJamku2DJQTh8
BEPweRAiOOnzsZWE8S4xSoVrl1Q/t+fBbsqKcLp0qfhCWTm1/Szx5DZ3fCM4nQ7zbiM281b8nLdP
WI3KVYey3D6DK0oB7VxI3F8jRRbcp5ZNOyq5Cbf2BgCvJ9rROjCL7KWCFgoRsw6+HgPElm8TNMDY
Q9WaphxXC1KA0CRXihxFUZng56MlL93RZWJdPLMJ3OJp7jSnVgALMIa4vaKZk3tjM9JrjUtbDN4B
I9nqMU0d1tCg3N6j+QCE2Je/qboZbpqsFfEjWE6eLFyU5LSJ+FLvMEycL9mOtTa9bUY2giA5frEf
NZE0WkZm1Kjwrkf8HVq/Bi3HqdRCnrGWnlSPahUJoi/zzpYiW7ijlsqYo6RQ7WHLPqIdDEeERdRJ
jV2HN2XpW1LwPXbai1PbXm938X4NdrNatI9mx1xGNgvOVrnZ9MITFDvbxEM5V/Azz1xQzWn18wXH
AJVjfyxoZ8plt9fAejVhS+GIIw7e3eKcN0F9KR2UUKK0YJfut1vTfVoBsgGCREHE6jZrDKOklPf7
YYjbPl5tIAixT4LrXLNLwuTXMLLEawvflzAvgY6ky6XyJ6fj1Gz6V7yY4XNQtniCPCx3lc5WqLuh
L5fyX4FiSlTWBH90+qpKWaFBtqDYkH9x9MJB2qwi2A4LtfavGcsVR9LfBdJDfdRJQNqeuIA8oBfj
Sm8UkPSW/dEvWlT7NLNBnC18cqqbC+2mOcr2FUDAYz+k0qGkdRHat/IiF7ImEPYbBhLPB3kSbqX3
l1HGOGg8XhmVDWyAIzd6Zz+qfwqznOneKNirXwvfK2OMDeqGgQB6f7DiAgziEY8+roryLfBxnYIV
igfnnwFH2OrnexU+jzW/q1Fx1OhvQ5ZjqXeRwz9C4sEFdgdozk/WZqmm5BXOXJAW0OQJC8X0HVDa
AQphNXK7cZ75MX0SwH25usduPU5UCd6zD5i9bcneuRQvwirKZj3z7QI5o/8yX5A/kHgWheKMVoJA
yh2VDIO9hr2OKOX+94660LtfhuO3MXYMzN2+cmqJG9uSfntD4qRYZh5gwT7KfoKNxshhGYeoPnKI
i30AJ1Vcg7FKU0oK2b4Q8d+Rd0Fd7drPVIyyCExgDCDzTM+1EENYXEl56PnoFKypz0dBrmEtgyiX
wIqXpIvDvQIllfWFvHZVZsusbwB4qFzQ0woiSY0NbuTUIaWoDao92vhpL3nIdY96VA2UKwBrhLJ4
rPmCKZroAt14gyLhjHQt3q15jJdXCzDZlo955nY34Xns1XEhV94ztm5/Lx3qa3x0on0nPib5NjqJ
qK+BcetR3lxNUGXAzLncFEJluPEpYuWd8kuv0uiyPkc35bUhXIXN4g7qzoTpaTLd8YCexMo4oxav
563FB96g9McvlRdoGNay9TVx6oqczd7+uYnbiEsvRxWegAdCaEC2XIUoGD2TPle54utfHgCLRP0P
TUlol69ErieksBSjkD4SCV2Troe7qNNz6VH23hrh2yWzZ0KtE0af8U6WZEWyzP6ZS00Ic+JPn3yT
Z7KvQlStNGEChPKXrVzkRzZwYCEy4wQq8R0PBEhiyi746bCX3SYkx3zinFXtnMEnLYSzNZHlsjyK
H6WyOXs3iCyGMOy4DIsL7ic7VYlGfhzBlhqsFYE9pCEsQJqOEen74ulFnDZLhX2iKt8mXOa31if5
dacibPz0oaWSrK7sqDkzFG5RfuNpNoGPZM4wzRX3dEp89KsaFn2dSs2BojDYoC55nR5ndOrQvHyO
99wAnWuUhzTKuKgg1RliW7HnNt1UKIMU7VUKN1q658wGPck5ppU6Kp9cK16QrCp/OK6IJJ4Up3k0
y6ZguPMnPd8UANsSlrafWw/lDklzz3x1yPQ97n2unXktA4IwDxITKEaG+cjuQOuqupJd0fF2LUZx
NgV9g+SFVsFtO9DmFLIk1337DrdJ0ZMWVW6JDT71Knk8KlLqzXaOU5JEuQaOK3p+XgW3bkAy/JI5
lmUQR0PIbMSwDkooA799iQOu/r0mKDf7Dx6ApX2OJ7nY5p+rUC2Dz23EzCnIOGog0fhK3D62q6YV
RvUG9j98hINkcvhlDogZh5o7TbSeeDPjSAfJ9Pwlv9Emh0Zuunvpbvs0lpeawl8IiXYhkdVBfxBO
hYdLdWFAbPZzsXNunk1lAutRTO67eR7bmkgA5qf3OhQtvnrgre8MQjg0T4GbT+mlwmpTbK+sx5Iu
0R5oUGzqaf2QTeKB0hEodbiGmyO6jra23mwdm9omx1u7o9X/BjMuc0mOq6fWLnHv5QVE0H/Tpgpz
KGTWrSlhLUI9cdXqg3y5xqeBjIfAto3jx2KL7ZSaXDXHinq/IU4OqbP3dNArWspIVBUS2TtcVXg1
3OFDE4IX7GsCexwHHTGE5DMFSshJpp5kS7ZUmdrH0t5jWOye3ZYR0ODGL+ppZbboa+rx9IgV2zo9
tya/9zmW7zMq/VrcHaiMCmLYEUimw0K+yyF7oz/T2ZE1RF1DhEDwJuvpD35vyPzv4j0giwiiuD3o
FSIzNWziaWQZ53hUAS0HNldLck484AN6OFZzdp/d7A6HoldQ3Ryqk2uwcvuzEA+2Mz+YLjrHmlvT
4WDSRx7NbhBN/Fc2v0x9JKUPNGowi0G9GxG+0PQcck6Vwn+4dvasbH6DnTLMMG/w7s15ZEEbTfau
wFM64OtlEqTY++NiBCchs+nZKMBjiVbsYMMOAvV7kz4aZaBsNu/yQFAK2Y8WuOhhbOmElZdGMnoJ
h9AenOvLQVYjHvKUFIUqUI4GG/8YwYYgp97rdLKsZdquDU21kKtq+Fk/EFFPMJW90557hTChUIUf
NDKXN3teoHYo0bSk+aM1jvAzxuufzUTCRTCO3bfIG826AntKlgKQCcJk9Ym+ljRMgLdNvtukFEn4
TyFGRT99QdSBdSxluNyWyJnT3GkkLWUQXlZTk89PBcStwWpMfkr0Y5ttn4TyXsDBcnyO0AyPe70/
52PeRnpXOlg9qJEI9Zu3iymtPf6Hq7CyOAI1OVq8SWsGNA7ix3IHnnu4EDa1UXi4FZ1dtpGBmcVl
rU7TtgOn/ijAho5+ZbsY1cb8915uUEit8Doh0OQJXiz0XTx8E8AMdvCrV9zcpXejBk/nkwoBsGsU
dblI5kbEGTa/QtZjVIpbS4/ZplSyhkRJH+eumG657dwPGkBHZHJMKAiPu16/0xjYMyL80a6GF6dy
uLA0m92p9bbJzocimChEhqPybyhBsYm0lmvBnvrXEJtrc4fgv/JSD1yXf/795FjK3uVUgsAecR+Z
20CVRAMemLq1ItQtLFLS4RqORJg9yi8uE5Lt+rw8TzLomjtgizDruAqiewUAOFOiYgCozXtZvh4i
EfszJQfoqJdPpppBilhCv4d2AqE1LJgAnTIAkLsquHl+Ydb+pviC+2TdmDmqJygs6OuBPqIM8oSd
plwcs8y8VDHKvYh5L0N7uhMyt/ttM8f2kTc2fzFnIakmFifZF5GoqV8GRlLNjrb+gze8hasZKuKZ
FbvD1WrqxC6STxJeMJT8/gn5osXmjF+R5QoD/Usvqx8u/83goZhwS8uACcJwAsaC+c1E+tlolPU3
zgKbWvZXQhwxddjgpowAhrWDQU64KWd0rAQZJgbuI0Of3aQ0PPiqoalO3STlBmgP9VbLcgEUCizn
gOHnZwxKPtHftqoleDF736r7x0J468h70Kh5JQwfvqMy2Hl7rXH+kovz1ReB8MhfreKvAlY4XrVR
sD6goGAenunKgmyQRO6UpVTWZErGXNa5J5Q9gDgMoKIAlkI5pLDvjUZZ2n78nLWvrRkw135R61vR
Uye9vW2CSAKYucque6GSMvYkjh3nwY54/0Q8PVjjc8tQ52ElmIQhgW4Acu+Na6G+DXRQ4PfWkhIe
HhvXLl4Q9MrDKSyJE6GtLpHySJktf/8TWvaZsflIoCLk6VBLoPIqyKn2bPnih+yXc1Slux/GgXCv
e2AueH3Iz0xnz7GD4vs9NFm9GGaggmvai1WGE9Q4q5W3fCPHkgumxybGnDSr00M3/UeR3gi0gg9S
1orBZVEXfxSIaq3zqdKDGsk1g9PJ6E8NcHGbst3abPZDfEj67XGxJsDXHoFhZxZjzbVgorEpqCei
miKzULBXHorQzRyGJJGJ9g9JFw5bAhXQG8dtjA9WoxSDAzGwxb+NogERCCV65pJjxiFaE8It51h8
qb8btFHiI6lqtYfu70ZscalTxS1jyXcmIHv50AsrnT4xLgcEzsDV0crZn685sN+1vpg2tKRXjuF/
gpGkagQuUlWYcTk4K0EmBbw9OC2UEp7BauJNHSBp1DFD/nlcYGqNCzM6EkufUxZGPFbdS/9g/pwM
6q0DZuW9BNsLYYGeKV8bfIuCIXuwujy6BjkQBX/1yq6D21A11fTHDdqSF3Cd7zpu4PJGXZnCry6W
W7FBluSyoVWB6UePtjogTt3kCrUnjBkLVDA0fTrdtQw/W2xzS4DOwOiRSPOEXt3CTuEK5E15nDKT
qgi3Vdu+ZxyGTZFeQAIWun5EJwHdHTrwfT5vkfNjZCmksrycD+4d9VusqFSQPnC7Kt72Pdmt7YZ5
4cYmrdjl7eJcNlB5+eGrzo6KpIn2WaCo1nCto8RsOKLbdMwIL1ZImkYo3DZvZULICd9DoI3/DEp3
JOr6M6VgtgdzyKo8+TQR3PIYTmBY6bgPkwQPohtmyhWuiFFQcpNGN2/Mb4maHNVN/Y2i84jd7oRY
ruh/yNJiy08hFNo7NynZ61BP8fniy5svve8mIJMQEd128JBYoYxO+rGzqrMQT7GCof6oL5dgZrC9
tRPM1shhG9P0ykxgSaHFzN5eV43A6kHxPeaUNvMs14tc5S0fClkWmOSCTcaN1fvjQU7oWkKF6Fe1
rNX5crMOdHdomQiLrNXr9bciDfwWS/IG6p23jY+6QZV5L1mtgAHALIMxZrOWmKGgSxXrRKJ0lIA1
DSBDIEjo8UuvogEmIPuUTEfhgUhVnB+Nzx8rIxI0vCI444CGtLxfCBIbIOlEeEUuwqpgnSTREP2s
6qj9UfodUmTgXdan+4uGfoRWXdm1F5e9Da+qV62KMB0jWuYXIoGCng0XPgIx5ITOP4Dw6rbLbpHu
vZmqbnyi4LH+wmyGGilc3LnESb9zM11O9IfhKVhU7VVUXSEPrdbZtYBw36/bSht6UZ9FxGAzlHym
B95vl3mXT3JRJM8AzTDRmWBnX2l1kH+dvitHFKV8QI05u5igoiLSyeaNkQ0LTz3UVtJWuu0nf/WC
FW0eb3J5lIY8+qRQ6EMp6HanJTe6RVLPoc/OhDU2PK44eSPuYC+W9N+50pcWJYwbWPR6ZhxK5vv/
Y4DtqGwiwo7qtWdg3uzDqgbOZNNGPse4khK9MrPwbhdN5CRg6/fjh7WxEeRtv5u3VRgYibZtZaaK
CXnv4Cyts2G4vjErmMnsOFPTTb0tgH1PF4UWSmtyXrmJYfrZ1K1SUBi80vQxjFzWQr8IUsfmFZHR
CRuIOVZMdF+FNIxGguak2GAvReyPA6DHCX6AYrFwgNkkXE67BhDVDwRq7WL9c8nChpUPepEb6Luf
WsWXqYVMCrM6mjx8uWbIkcw/UF9MjJUZEPPuT6MzAZ8A1TeTQVu1d6WLId2IMqndjIeo65PMLCNU
rxQJqqXlx5W8A5/UTo+CXclOu4qrFOsHSsi1qWaJY93t5GokD0I3t0nbobw8+oqMHhXOX1TkIOk5
/Tb7gYhI9jiB02KVsCeOc8lpYA2jEOYxYJcQ5NXPfaJHgcZTZfO+CUa2OhAHc2aD82oxjKTSQ0lW
LtXeloLTEEwkaaeR+Td5ojCyurktQuqz6RcDzk25PLdo3vl3n6o61wSqEHfUzxtX5Q6S3HdZ6MXP
jUoL9mIDp2m9+OUrOS0rH96iWZKMttciCznaRCjp93PxI8UukrJ7jp6/vszdgrMNy55Qa3DBDPMM
+FUN1OqLGZwbJ7UEmW7VGy8Kf8+5NNepzoAXVKgSc+z4RTVGXeTkWnqLRjp6/IlUr6TgcdvKRxQo
rQYET4Iy5M9hGkULBIlr0N/1ImMQR80FxGcm1kHb7TZnO9P9gPASLCqrvSFmFQmCip+dL+abIOw7
RINKZb8KX6t2KSRz5sgRJtHdGFMMQGFKa8tpIzkWhL1Lj/zRQuqaLdFg9T3AJqiuSVOmp8SPsKSk
zkLetiH/qAoBNQPbQRSwCPvVJqLyWaX2ER+B4me2nX9BYl+DXdk/JOZKK0OMOf/+snwiNqHKsuMX
D2SobBB6Yt8z8o7qVKHMeuJgoccPmkKUX3zfWV5RcIHuUi1FmzQX7sm3+hL5QcXMW3LjV+8hAz7/
qkQ3zs5O+htboJUJqUHxB84444gKlqyFX3Q+VOhnSI6nRQD+6/VVOLGg9Nd7WEeNx2uQIM9wySEQ
sPVpfkLpWdGTZK9OIJNIH1aJYR3om7oDeFioFi8MmGNI6pBYqtUl3MXf0nrmykRtOY2h4wX43+Ew
nz+f+hIn5261pA4d0f7V+6nT7wQ/+LAsAgJE6RgiO0lO0oMvXz5pVHGt4uPFzp3G2qSmSD6smcl5
qduS0Pvoq1uB/jBHXGhhzZePMlMnCkUhY53XMiFMU8gu5Wbg/AL1Hl0zOdh+uqU7h/dtteiqwuzc
kghRR57cqti9yAWM6ljMHAaWlbCufsOebtynHNNFYAoJ3M+TJ8JQR66SXWHdS33Yt1xIYOMU4Y2u
sDz2cWpyNPjOOc4aR/GF8lZzFAiZd8O7a3lL/B2uhekU3N783kyG39JhsAisxl8hLCK1AKXr6tdp
B6CwqG6+TqPP7C1y6ZG9bbroOfcNGPsmxTDUUXj52/8WEcyKpLLEAzNfr25fq4L2YVzUMHTmV48y
jt9tIgRpfjEz+UKC3bhgUxyBl35u66ul4UJedP0Zmn7snx1yC5o+tJvbmONoKnOC00N1dA7nFG9C
pWspktYskBzuZS5vk7/duNibnnbLQIL0aBjajNdBr9WQSphcYMROako34ELflJX+ayXRUEzZSvXv
O7wSZQcMV3tGd4yU5KjumzEd2jhwhrs85OCqzVH9MurWfiy/UltbvBoWlNbGMNSrobiaBKf9mgYW
1wbCeAhkyk66pz4om8G8zsZP3Lwir6SPdvT28YAotl315xCmePJQNKNlJwk/DuKEP/8Vu84lBW8a
7zqQI1wIUnOiyb1Of4W6YJeeOZcXZlglCLUSmDXNTve2ewoR28Z1X6BQwMuk8x/WfSe3crcA31ro
yX20JPq/j0jXXb03ne0HvaH1OmLKFjF3BIzE1jC08miWxzu8sBAOZ07guxVDYa/iU37WYv/Pnp4O
scDo0ZzKqln4gIzBNKNR5nZzW+r8UAJednfqZu+j1kg41wcuuyu6VCOEejfmkxHUtS9Eknx93EEh
iqP88/+j6CE8siO5bT+ZC+r09+i3Wx4t3aryWTAKEp58QO3qzcjgsLMVdBM/DaItzLpVXLefZLPE
yzE87xR6iAr4C7h8zN2bPomb8e9W2OzyZc3GAYBKYUsvvXSGC0TskcOWDFqftBbD+SqqtKMCKsTJ
ywiz7rnV/BXXwIIcpxqz5Bb7b+KcbkxPrAxnDP5gFGy6JOMQScVDpgFZwnWuqunqLFPOt90QY/bH
RgLlbCYHQwYpggdGdNHTKt0mGxn4kH4EJr7WKfiTgI6vfZjoekjCD7H0QPFz95xTKVBX/h1MWxME
KNVoN4OfPcslO3HfPVexPq1GPEQQX4kAyhLtzH+VSZUVo94BTwh0IOqTkHaAz0sSUtw9uALZgUHp
5bXI+hIrF1vV9Fw1bo+kH3JN5cX0mglzMEI1HtkIVPqLbUbhGzv2cmto+OcQzdOwOPH0o2I4Q95v
Fjb0CXAWvHB7muvaAxrn5JFcpCSi6VSGKBl5LHRA4WiC1+easE6zbwNpZxXeglaFKwVWD821M/Kq
Mj3ngYl3CHAHgqrSMwldDe15wjbYp3BqFLjoBmkjp1sTwe7vkFi6R70Fox26FToMN7obfsaQolj9
B+WhTwLSir86Y2Q4idYD/8qt+hF2tvx1a/xiK7fYJFdkPJMqopdkKygC7Mb83QTs9PPdo3NIXMH+
uKwKEzTrgA0v21myIOaDkl3Cok/2gpv8+fmp+PQ+ZftHxXCDjcC5W0UTnmJj/V3BoK/EOSWj7NrQ
TR0/JHmjQXJHv7zE6TjKak8jmM2d+9Jy6KKh+SPMljQczDvNZfZvj3vE4lR2nNw3Jc1gjAQWZMjk
6PwMWGFdVVWeKE9j4+KZQPcLkdmWkqCI0oGis0kduiJawuXABgvU0rLQqjTwj+1nBi1yllPGlVCJ
p+bPBaiBBji1ph+TUVQxb9LDNA4LKjRXDADf+TMZMiaCrDybhShBq/+vdqvXwGGUOk9RH7Xd7wF1
I2b5/gNGBbjaXCBtFq3IspK5LyA0bgx9cXiUIKgrssB8PiI8eZTNgW8woJhpA3E0LnzXjKZUW0Yh
7LmZrYnHx97veSzrDVhtTj6sWhoavlkzQn1JaOaZVBUEatZXg1uSIE/HLplPoNrz1RIGZ4eMWnKO
rHKeUw+s+M8cJNPbxJ8IbWDWCYW4G/sO47CoJeBEnzHdOIn8AQnR7G2KY77terPl9Gg0ROOwrUuM
xWBCzOaTnD1ThrIaByCdn3SFWHIiFP6Pr1Miyb7iCpKeifsvv+RrVdvTw/u8C+SihafyC7kCAWJ0
MVr5gPfESONMPzIPTGDT/sH6btQi5vpHs+0vgdKzkqkFn25hgqxvD81ZDigS1002M5iQO3DrXztQ
yvq0Y28PyCFSUwQ6GbUN5gj5Ugc99zuZjRsBRBk+YAiy9CdRJcL5Rn0yNgl+bgF8Kz5zDEwJ2W9W
iDUVpmnd4s9BVBtDbYWco0hjVQDD1b7UK4lplNyL0jxt6o7VSZyzP79AymB1h84V1vo5UKNS1jhV
ADcluShC9IvQhG4P61eS+lWCaIS2odTCq9sJ0FjUlKjRzWhjmxlJLQaUHxxKvwLfjzDlRe5CvgP1
VP3ekoXxCj77E6pPvenz4VU9kVFKEBquKYCSCBnk9vmCbPJFu/IUna50fEO76VCW3Lux01B4vl9C
bWT4P5jgBGBMsadcz5VdhdkcAo5/vawwgAUjEpFH319H45zU2AUyJQjCtK+tOk9tiQm0Qx1rzT7R
f12ZvIE+gFSTVlwltEgaW1d4ePQ6aWGJCxifbJzOwhXc88KPfeTNSX6J968CVjTH6KA7J0Rjimlg
jG58kBZRCOxhfYeqLB6SLh3bcGEH/ePTyYYLj4OnzVGW6I7GyhN77OGT9gQ2OxTWWxhgsGAYHRQQ
oFZ8FFDZR8uZwzOO8lh2gZLBNYQ099xjl/iIFtCfHuFM3inpzMoW1XJ7yIwCal0KfL+Fy8s0PjGX
m+C3BVh34EZy1kSMpq6fa9Pt1uMhTWzVAgtEjdtdQv4tlN/ymPjCSiVtpX3wqiNH5nDZNAuHk1Iw
PPms+un8/qMqQLwvdIccCQ5y4obS8bQjfwnB30MOEVNSirC9xcUoe+OlNpL4gwwTcmu8KpSDKmtf
ViWHZFOCQK6LqpT9PQmo1VIcTALUPx5GUWGFuvGrHNh17vLWF9qnjfyNJFO3hHLwGCfzJ0kASXy/
xBC6i/D1qm7+MqwENfm5vJgdfQMKu4Gd59hzDFOKQNsTEXdp7OXaZHd1PkHkWC6uqQ7XxuhOrukK
wgbowJYY8uXcfvSq0T8PlfJ12D5xpVgEx2Li1YHCY3H3I/L5lRGqoSSCoS3SsWEb1JrcDP4D77up
H5s2uAtx2BEI2FqK1OjiX7dIExxrj/U/YNyqLEtfxB4Xwt5Llc+dOatkNqW/tG9JE30NxqSs+XTc
GSllMqZDHRLIR9m3wT+P9dS9gLn/AIAmY/KjJIKf/3dmZ18z7rQu9Ad27zBq9+WyCLMwoVx8w+ln
WwZvmXtOO0Idh+R9Rd1CJgiWs1FSo2L47LujXtp9qgWtig0P8fPoRnfqLXgEoTZhmV/Ww817BR1t
z518HkkCiroRMdm12kp4pbPEUfsQX9U8P1e4NDrYBkA0BtE61HjnuJwEEKYARE23LJwK3yzM9xl/
JbjErjoRe37AaGKntAfxtb5iNk8skbtBPyu85MIFdXwT/tbvEoqNRwgcJqj4r0GP7LwHSwyej1GA
9an0//Y82GBZBW+2rSttwsPNuyhyHFKMPw/Gzr0JVGi2a5jQ8FzAtYDYZ1nXwhyaiCMeeWYs1hFq
FjIt8amCprMyQ4fXQ4V1W29GFR8fYwx3d+eEu9C9LBsGSU+9mE0P2jJvsI7fuOywMl+FT3tMf/p/
u7EpV/8LBudDTzS86QP7Adeg/ZT3Be++cKx2kvSJq45gcxn5K9zQOVegQkV7oqQFtwsNWYiSpS9M
7WoNn4MIt7pxijNc/WhZcvl/XtkPa3g82eFQIoXWXAgE7CzZ5AINeLPvXS40xuJDadhq+di81JBf
9GCazsd57kVPq402wTdlH5tr0mC7C30JrO52oVA43pnulCM8im5pmFW0aeQMjMAyTObqmtWww2HX
saAOLvDkamPv/3KlkcdzLG1MwvsJxZKlCjxO0vunaRRFwBwcvMRX9/oh376WwMiNSbOGdVXOBAGS
K7fDHUjQDOa1esJ+hdtbxjRvqzIoDbkxtYRGDLFLkjEU9wUs4+yov+j1AQH/QXeOs/XY+nFpYnbg
vM9sQWTmbgMKRiIgScmEGl+CZD8DBb6Jx3nTpJrFBPSkkbIToB0cCEx04yEkZ1S99jEhzYTi/uIc
9xCgw/sBb8L96YWaIn4G020KG02+BHbnCvnNcrf8dXT/qHuUmeDkPbMp+tpS4si8WwhhC1vQhTqg
OPd9JbJiFIkvLnuYTVB6ys9rP/M9GDdOeRoUo1UrqL/LU1z9XW4VhcCpKGEKEAnFjTKoABYxddwT
9vSihb64qZ4bj6uhr3rOfZQ45xMebXvm1KRT3DGYv1aA61OjYK+tEZVeqnfxWUVVgoifRmHKVGbd
YqrS2Df07rMZblqc93g0irpxBnViafDEckAa4oFjPm5BPUySl9JTySc/BmM+HD5Jd6BRmGkzfSpb
gs5hAIGSIXkoNVzMHcJHCkI932fdkcbPY2HKmN6mKLbmzHPSjz0zX2h+80hR9XnLKnR0qqmvrAg+
Z1+6Gwq3KvwBojkRiEQU6QYbhjpf4/pIzGxzW8f4+inszViZt2h3RXD6o6I5zUSCdCZgo8XZPVoU
bKZKgqun7kE9ujW6QLp6iZYFgoEMMLLCpFjtjAgcIB+ypX1E1ZmM8AzB546CNyQlny7yhcGa400t
I837yTtOAM3xMb3KSzD6doDxzVofdAfCPN3NV2tzQoH5ef+amvoW/kgEndr04d5N/S/3Y1fAZ15O
f+YJtIFO9/irJTeZvq2AqoX/magdoae/OiMg57pVw4o7xapAQSi3bHSqVbfjdo9pH2l39fqzFASt
efudhRYe+hbDxXpcCBya0eDm+OHdjCv4p9OrQt0B8ZoSpqGwX1OTLUI3tLog4IR41rv7pBxpDtkk
vfImPSJIpWSPO+l33/2rEG9QohXfgp740Nw+IDTv1vSzJsJs8Jt7OqBCsBOD4BEnLW5lxVm8GVUp
WYGrKnew3MmN6CatCA0sk30b3YkR1eFjfBXNAKAcYbDgICyAKlXFueGr/+4Z5jJdV3+S9TEIU6HN
lGt97KKkmbgrCT7xrVkWJ5VDfoUxDnBR2h+gV8ymVuOtRkweV2RsjMbDpkg7CqT/K6blhjlM33qp
Utb5XA9FXPFPqw58KH4ZWkj6Pg3ZddTuBbus4qVFpygjB4h/uoIVk5hee9HHQVGvD7QDs3tls/Qg
BVZufZXWAVCCLI4tGCKfElyJ7x6Gum18A/31pS1nZNv9dEu2kNpeSNO1LKEOT7h/JlqhSLcqYEKN
zXdksWJ+on7iGTLkYasB0lc3mnVjaMiCPfp4PbMzm5lCwYh2BRZSE7Sqcp4gvVWgMl5CV609Kkt+
+bLzNldrR5pJxmqe+h8R94dX1dcywfMSqROemh1x9fy5ZS/PD6aGlqL5PLqx5SXTtNw8AXXs+fFb
aWCXCFr9Dr5RVEpdnet4QJmshDB6tT1EWW4PXzUFJqXqit1pNBGKkAH6svCtV6TAYCX9T22UIfRH
xFjfE8bCOZG0jtCR4N6nMfO40g5/nLOk7nvXbiS91YyLfDA23gPlII2gJFR4tMWnzQkKIU0+bn0Y
omthXtT+1RGacSSl9uDbkQVnLC9cSDog4PRNMOHZypz0Qp+XfJ49v4jYy7MZylvqC4qTQ9Dqhu8D
sglg73D5a7P6hWYJxbAB5edRrhCuTqA6UzjU7dG4PTiKNKu7J5TeZHHVI08QUykioN1rTSXBdESe
k0NF2jZUqp7jWKFnsh0X0DimQaHbFwAl0fZ+nm0UH9/nPqdDb6Tv74s8qtK1AI5u7AkgoXgE5IMx
2lozL6znpUTfo2f+C9lRLqrGWUqBsXeAtZEdevDJsDlKDewLhSR3OFPsK3zXJpLwjiDbWHB9Jgl8
HaYzZ5NUjmGqCyt442hXNxbanGTyXJ54UOwWja5w2ZKoBdSkn0h/aOntF9XM6Lt7I1wXpaaOYx9T
7S6VCo4CkcAPSQu5Ar08eUy4UvnyjzkY757OBbRBSegMDuzChqlBkl5Ta74uAl1G7S/9WOfygODg
RQjyrnUwffv3aPw1ScoxwyS3shqaf0dSfE8vwp1Z8T2no5TUzRoXiCEeGAGpiMODlqccZNh63Om+
83kQ10B4xe8v+WdmCgjczYmRwALwk7Q5x8FLVR46r+wTBWQB4eMNAP97dVy//NL63FTOL3LZ/Kvh
0eERUlAslPeS47vU5VwknZmwAk8ta/18j4sEwtDklHKsheKFm7UbPnEF3IxaeYxNP74BiWxNGrtB
rdLxQ95L5VVM6ph/W63thJLrwDEkUBXatrKVwvaiNCS68QQZ2l3+Qs1PWgd3Hddw1o7/of1nB5UI
8mV2mtoi+Cp4GNcOYm0rK0D3FHDakzGTkcQrIPYvRFhxqjgsDu2VqCT51qeTOZyG26PZGbJgrGMY
RPTtHPVXAn2N3OrN0dDXMvti7dxcx7gDMkumSOodSVg1/BOj4FD2MnLELm1QMZCXNxsFyz6iZnRV
4h+X7P7I7aI9d0Tq0RhmoZPFwKA0ILy5LBa7O72K+tk6H8ekbKncSw8/gbaJUkwR4gNnb7cd19Ng
VoxmLayJY3sXXOcnoAVOR4oIw1WMAPq/ukmTl8JNhjCun26Giw6ChKShqF3iN4z/Zrgcwqa691nB
xb6VtOcLgltD/CgAkObrH/Km5AgOAD+xCUqZzHLD3h7Kg/9XvBXfbAa+HbezFOVYugHTQLRSrCvp
Wg93mTLjw7TRDd7xxGfDKfPhq6nPNGU1pnI8l3rFvKJKEjN07ztQbpV0d/aGTqgxHtWtpepONIjh
UXIAGY4bgNLSb2eRikNxmeazewqW2ZWbHielB0/V/qwIRJP/kOGXCJPZGHiXfQAMbEh7FrGOXnKJ
mqRQ0+I48hDRSyNU4GpwvsFWc9HSNXaGLnGrxiismca+/6OZQTQecJr6NXa4vhYDm9h7sOdZbcW8
QcbYJEp78Xqy3OJO+zjhKzziBm2nAwyk5LTM1sEZq9L8Vq2ZiUKrY03lOEYSJFq07Bt0YgGQzzx5
dCC8UvERLhcvR9PpmagvPzk+SH+zEYPyZLeDbAKzHZJnpeFcRqMRilyXgkh5tMcjAYt6una8cIzz
1BzyO90JRWWfmYg4hpeUm14yesNtHiJcxSjnzaNAOSREh8/l3pPrDOFNDaoSIJ9UR5DGClPiGGvP
0whZCAct3gEF36M7wQGN6l+kJro6gv643ygWZxIGkfFGW6YVMfPV17cuwkzX5cQ8Pyp5PBf/ZA8L
ebMG9Bk/MLiWldUWeqzk/RN8BusjaP6VMaM3LbD51wk0P22Jir/gzyjcMQ2gBNxlqru4hyznp0w9
HYFv8ouV+1l7tiZlJAVNvXzmA+hfDMP9mA3WB++EAL0+/CISDBQLku+ioxMBN8hqd8OhiTEcOowo
UBAEf8fLnTOKSBPk2il92vobQhEY0qiEdEVoU0Pl7S0tNNcowTHQIBQNMlESdG4loe9AoiJ5s2mY
LQdY4NrhlvbOogmYEXoRuXPc1yV/Q2e0+km3Fi2jdIk4SuF7LF5cSUVc6jvNCjEZDIgPspqDSVXr
WTU8ubSNbejx8LByf8Jxk8NH2ZligJTLtpwA8Con6i2bg16PpXYoFe6KpVBy7CrFjinAyyglKGac
hyTci1F3sV6d80QrbUD0zMwl9UtOoM1Ihp8u9I9uWXyu00/PksYQow1mKO2E8CvRZwStjBrn95Qa
UOHUo/HVn4skJiZD7YmjgwcSb8sJy7oVSAPlJunw1nr0aFlXvWCFsB7jTlFu1HX0xkKFejCbmOg6
ytVBJTElX7GpcFrwx/tKywgXx4fYQ2kVZT/njHFac0f15IVcAtqpXMuvvfP/2QNBxDmWo+/pXsN3
rJuHrX08PZ16WQLcvUsSKlaVDa3CHfH3cFZrweraWf5T5UI4+QOarAc31n7k/34njmq/1efdZ0zM
3JJrqVJbHlYs4VRMJZJTt6AvI5qLbwQtZPQPEHxqbqs4/JWBVtmJMmDuDcptWgganB9hKfpqzVaO
13PH0Puerr/SRvkt8cuTfEidhXjRdtN3JqyqjszDZSfOO89UhiM1stB377J5CSOItVEWrMbRovVX
T5968/FHOnrLiHaApbK0GFwSJqMNuyp+V5vp7qDN3G6Uc4i1Teq5pozegMmnf65eeMd6M8dp2/IA
nyqGbNp70LFC9RR0g8mfzhMPO8TvCkMWbRjvjzhjALVA9CcGgTTLH09CEPUj6XnbAEm1O2hpyoyF
qSvPYt91aHNf9+NqGzJ75ROzUbw5RnHm4ZjLDoVL6hvCUOkLl0Ypsm9SzbCdC0Jgbiq4ZIJZkekF
Rb0iCdDVyIzszyISU9Sq9nZzgruv1zQJ8Dyno2/gbFbDQjxSY780eG5ydMY7XFDJAPI3Tx/rdhQX
bz0qrtfyQldRMlHus+YyLPJLJOMlsIg0NAhS3gY4dfBB2Z5lTY3WLIA1WwEhI+S08YDRHNksiZxA
IH1/zRJhivBfKGxjLxP/z7mrozjrhroNlfj6obOCPotn8gCaHMs15Lr17JJP2+SRgETUtayZh+d6
fsOZttdnO+HklHd2K4QgR6tFOCmwe9uvy/6YMdexGLJTdihCl3NjScihOEuZjVZUhHu6v+GSGL1P
0GA97GDdDD6dRikoAlJk3haYwFh+V3ZYykzYbr3Jk/Vo0rNrEUJbZF6aEnbr9EAqP85QU6a5e575
+7j66o0jobOyivXh3aZHSJ0YsW83Fg4Kcs3mLGUKeh8mwBMdAz6Smcd2CmmJ6dFXTXOZMvuHNydC
l0x9Nb9uCLdxyt8gGm0rmcP2Gj15af9wDEy6IkLa0jBRXGAuFBX2C1cTfGTCDiMx3aleOYvXeNCT
MCv6t31gCxuzqLCQjieWt0kknw4GOm8s+z5yJ8B8CuZgM2pOh+ucLkGIw7ZuOvKyGNtTEsMuhOJl
vEWVYCxkuoO4oijvwxSjEHcKKnkXrE0AvRazivKb074Zhz2skrrCx9hOiLnZds5V5lNgcogUXmcr
gfehESb8m6bmVp8DiYriIdL9ngKBV2xQRHJ5Hs4zkJPzd3t5nd1WS8PHLjx/rS1rnrAFVBNDTBsq
HDqHWKk9003U1rRLcD0HzGbDfYbNdByRB1jbRfZ3T3vHajLDAv68R1UvKSgcA+/1abU+pZ7JKrHc
5zK0+X+qpL1q9Kc/QBNQDN9p4WHKVdQc3GFjfoYlIO4fTptr+ruizhW2S/G4ykH3X7Ro9FWjuUsH
Ji5nk5k/yXVuAoLWTtIcD8lsRd8jaC8iFNzzO7JkLKg+htc5qQIUjHpUa9HTABfz1Xcu2x9P34bq
7vHCnN0aO7KjMpy1Wx2ZEvk/tdIuWBJJ6Y0UPPVK9Nu5YLpsEYXm3DKSF78FL6qw2YwicFShKq+F
nirxTmZGs8wAJTyAJ1Es4uCqHtT+cEizOxiaope03f9IZP5KX9Kg5Qh2FHznkBWTy70wyw93lG/d
efVc/aGVK7UKFKl/zISITnJRTUCvz5khgk1eiFImzdCvDd9iNAlSdhIKE8FhZHXgOqJNtnJcHwSd
ZNyFXAYAk7UHx0y9xj5lJS3WdIF8PoAWT8GOdCS8c2hiAJp4SWUE9vYddWuqaQGLx941Fc6JYre5
q9HBTpdryYzSt9KVqfKO/YTn5vVMNYLH8qMVV1oPNTkENJooQjg0KuhYOvGDZk3zF7CsdSqT3VcA
bbewuF41r+sSxtT355eDkYGLm74wIaI/GJcy6yxUvvRSwZE4w9JAP7iIjBdcapriDEaOZuEVWIll
TpsKlH55mnkEAiThH/URqIdmUuDmzLv/b/OyMY7VS+lQU5gXz5Cy0ne78PE0fn5sPyqEWPs51EH9
c884gjxcSgOFHRGBPKNsavz5wv+9SBSr/tE7JCyONY+5XdAucWlLTX2gbEgbZFmqRE01Xt7C0Gak
abu4hKlGPp15MvpjpYRxkiWnwzikaAR5EeQT1/LvXIctv7v4M1rtRucYxMG69q6WXaP8BxshDnW/
p8HMFg5okwp5vQMWeV+903ixu7XtQO0Imo0ytCUzDtOgRVgQvu7gb2r0fBI83uxwWr/T09uW5SXz
xitg8HiPOIjtUMQnhKOdoYsueX9LVjrWna/mWJutKFVuaeu2C1gch+c2jItIVF6kWGwzMcPOtRjC
vFLZMYMN1k5/rMcznETDLtJ7vIxb5cMxDpGr1F7FQkp0epzg927JFWuuqk+ocMCdufS8sP2+kWPr
cpE8eP33hcXJS6aQtTKu0lNNiZKgzz68fwU0CUbCB5Mfcx2hE/eF34zRX80C2LzfBLDU/kEJuDC6
wbcf0t1Q/5vIkKXHgmUkK8gljGUVOdahmE2OYglwaMSxaxwibBtA6bqKcbh/mo+c/81VepkOuX8m
sCdhKFeUvINX0SvI8ZANDgs0WAm5MaqIxnzaY27FlBl3AVOP2qPKIsbBExNdqEKpWKL46/6ACU5z
UVcgzkhR/2z4kXlXLnzkyKYLEVGTkfJ+OkwgPX4mZWI6levQ89J9uGOwuwPdBgfe+Vmqi1WAgPsJ
muikbMqs93i08MVlMgi6Ch7CwPtAzBJRUWyq5S+iaIlYGdErcGZNgCunRhUSKAzx3hJmSiCThD5v
AKMSwpbX2e5Ndz7araKEMpPxSqnaa9g+TZxpRJrnUAa3Iddp9ia6XaWsRlLkXUyfSe10iAz2auVR
JDInqm9kN1CW8CYHLy72gvBgjRnTd3qohY9s/OeyXI8PlfIen3XJbdXC9xq+dVfJJhdmcULmWQyS
jVJ/p14bCQkK6ZsxM4rTZOVVd09A7vNSh89/T7KuMqenFGvzXpJdr8uhNl77fiXAqUSuG9K839sZ
218YJ8EW6TU8FRGxFGw05jr6/cvK8eMCmy5INtQOOuxkSery3ncEBPaSEQTFDhaCAPglsqhgCqLv
StJoB63LxeryQ2kt4UBtvPvEdJ1liBwovo0oVXrYaTtrjfVPSUpsDtC28oaISlQcnpz7VY0TegHa
AkqmL/7PWPem2W5GDvbPrAaYdg83JGpJ/s1uz+k+t+Fd2ZVHFmYvnUUH/KzXAz78gUa6OVssvEnC
vXAwqTwJQ6PE70nKtvHmM+J7h3drL5kxlXjMnLvFp8ic74qV+4jwqv9uPXJh8g9qWTML1j+6yaSF
CfDWv92Y4IaSeYkoxaFM2+3A8nk/5HZ4+Hr82sWuDaBMwR1LOfZZwD/J56oHfUKA9TGmefye3inW
Rs653qnL/cPRf/qou70H7NVWLU8QWZMroa03eNUtZxbGHexUY+TrbM6/icRkz3MK/H9usJMslE9Z
J5THXYYKfhdhmYUZNIK86OQUAbVzuglRWkgRXvXRidmdGOWUcT6lA61vrlabvhHVSH3I+3JK9f7A
f5OPpEe/D0RyWryTdmksZNO2/uDzRux5x3segJ19RUmefsPfi2TzZyUkai9fAY1QIrXmvTxi8ew5
4Jos+3M0OAbFSEJnz6Nhcy7LIIp/rHK3x7cH30WblkcIGb87zCdMp/RpIsogANNlryjMws0Efro9
pPqeAOV40Ob8sZl+v3p/ZetFUhzCTCC2lEWOdnjUc+h63q/6oBa2Qyba51ZbxYVchiwSCReJWxyE
ft4g4TglJG5F+Ob+PCOEba1+Qth9+RBQWAoa7s10nP6Rcszg/LL64gpnlP4piaJ0kLLfs0C5ECRo
SM6VqRGW0cS0MC3Y4kdBiU7WMwJyLjLeYXYE7KRyV5nF7b+qJeDrVRi5yyQDpDCXj/aTCxVzEuyu
L1MtBZYlVqK05t4BESP0i6HtP+W8OLpSpULVP/DQzvPRv2l3nZCp3XvLkU18w+hyb/GDzwGupJIm
z7dKXvNJZcpI86ibmtgFd74f7h17EYqKyRUIelwrNm/YuVG0PVuJR193xxxhT6jE2AUSCRko0Odt
RBpE+XihMiv2G55TaPf9g8J+M2lFwpdYNf3PVus0TbFITxMbZTC0oizhqVxc83efdBakSbBfA4wn
5fZuprzK0A4XJSW0ehaKPPuzfgLiaF9G3S+GYnyQbhQ9Bl7fRGYxW7yewNbTLcjTILZucwuTagAn
Mzw5GsWneUbpVc4cpuodmTvKfbtTT0cbmixF74PdoH9nihVDWMaVMgNCC9WtMKM9XKACN53qFxKj
/VMyXTIny/m8nKH+oMg0zKljDJ4V55UTg6LdkKLVwb+kjoEvoEv2I042HxQRnRaBpWBrB984llgT
/XUDHgERYroYjf+3WAcmG7oI7M0N70c1Yi6K9w0Zz1wMLmec27Xa20lcJ8AMcrjTtw5FM2e6ArU+
Lgxd96POW3SMKDFrFtc6pqk0dlrI+4aSc3Ev619qT/i1x4FwEkK2lb0cbg0YGmFtcBmhRt833MYu
qWOgxWSZmRgb1qq9IQFmry2MV6YP4n0h62rD2J51J8wUpY707TPV+ACRe1LGKUp/r1xWuxW1WB3f
75BzQABxZZySj0HBEYPEII8qWqx+KjhDj3E8KLi7ntVqoffEC4T0+/eGjxxkrSjCYzJkrGkrlQk0
Gx6w8KP8+vEIeGF0znJC+zbkwelmcDxeCHxE1wKmbYVwenI4LRyasF720y94AjUYzzbZC6OvjA7T
PChj0W04cG8hhRK09alHUa69lHWMSJjYlANFJoSiNZu+6FHX0BISeno/XKZgWn+zJQa9Rg2G0fhq
e01V96EKgp5eT5BWlwWAGQeqefO578rG6kHcEvyLs56vtqK8416/Mmvq62qA/4EeFkAfgDGS/EUD
BOLEzUP1AC0a+opaRcrtmac0mm/O4wVsgKjqpsAMCQkZruSeQV5SWw0TaoNII1kyz8kBDe/V4hrS
krasGt7ACe+y8t4ea5xpUSrPosQobWg+Puwtr3QWulnqH9DUtt3L797KtQTT+XhvAfoItWCtYoIQ
KGjKlmgonTMgRezudfEiargzvEmL1zTKyEYoLMR6iTG6yorAniyu4iEox8m9/P7LTCksRirF+fTm
y+XX2FmsEl7OnnrPxS7oKWyo0ePztk1D2yiwvgpc8FuHfLizMvUYTOYKS8TLHJvtYenMas8rkUde
+MDyFA5VTcpjy3hG0qD1nXwDjjoXhi4AydKWTAlTTXH/KJrGrkYidZ6VnnmmwA8kKLdzHaiHOET9
/cV+nKmq1qfPwwyQWtNDKeUkRey8AWSvBXnWTG29EZtpTHNxAD9/HSXvbRsPUr7IsX4CtG+uFB9p
sOZCZ9OSPdsLjjqgawTwYGYGyAoCj29K4+lkrPhPk/uPHMUkhB4YuN2+Ik1O0rbDBXARTmu1h65Q
kf/vqfIRG2wgg+IMqomjs65KKhfxq0OovIJv5i9fsI7tqb/y27x1x2TUmoVEa9CVuxngJOfqVGvs
ADgw+zkoIUO2ud5u3pZ4VA6tCUwsdokQZeHVfGtWaPSUd0jBCv8DC/tX9kSkS+9ajg12h4hbZWAk
yU884BH75ZPsxE90OvkXY2C4GzhTCOkkaEKAGMBSjX8/aQAjATKA5RaCzJtnH92WjoWmOIHlSNSw
YlIOHhgpu1Mzwb+uADR8l5lM5lTPALCbvUPXnYc/3QTk/NaQQPh+rVbd9eRcedJfh10Q8z0eHw6A
NnZqFFA7x4jltJtZ7wFKrW1IJkw2m0Zyu0e41iNbE5VFeg/QQxFyWYbnHTo6FNjldlKW+wxVdapW
0jElGtcyuW406ZZBO6JhyMJMMLJQ/e80WVp97vQpjOo/EWOcTMl+JZjefnvdhknBGJWiMbuGE/qv
5/CNLMYwoO5QTFX0L25qZPyt/8VcqdKCHEk4W+4tU0WFjX14l+OnDR0/hS4rvJdUSF96FH+lNpZB
3CaQfa3DGtnMJA8kxPSCWNilZN+xF2OSDJFjOr5VNHRL+IXqcVzi4QEer/hIUPgCv8aLSd9Fohgz
yItrJwQx5OtN3hpN0sJGvGuJ6Caqp105fY7LJR7xLeHF7u98H+b3yD4u0R/VGUibrs2hqmsVbzKl
mBOFl7adepeuxMjFdOcCLj+G3LYvHVT5bhdu1dMG2rfxK3clLXTPykQYZuADewzbaGQwLBmQ8rlN
ZpTX9KZy4GuR0zGHWwEiiEV7iYtkk4dWNQRhuCoeZUA0akTGNbtGIUWZz8ZmXlhXunYxi23WVGlu
6ACMDkFW/IUqzC3XdU7vXwJ7zxG9+mmfLm1Nyc5Mmd5s0Ntu8cTOerTyUUyQ7YS4eUvzfuS0QOG6
k9vvlpanTwUGGUuGTpHtd+t8b7mf0TKmI6vOsaODP6P/AWaRhXGDXVfSGPKT+Giwlp2hlU+VdLPR
W+e51iPm/hgqJlxOcwUhFcl1lwSz4PC51MT+tKbVVb5U3u5MsJJqcFAgwF8cJA+DSbfdNETRH9RL
birQEHjeRDbTMN6hHk3k4wIhgZF6Spope3GwdkA2JwGXiA5XmPnWLjTpixo+qVPlQrdJJWxptxrY
wUUJZGVdWDUiZRDG6063RutO7yG56bv+9vksdfC59hBD94Z6iO5ov9D4b9lRd8k6Wq5XEn0MlQKm
EgkUW1/LYcdOkAx7vvOHzb6oZ06odP1GXnjeyMB4RjwV9+twPn2e6usMC9iKpbYXrbs9aBpPzxS1
DS34zD+RGdKtB8bG+PcQ/rRHHT+ee4pMJQmuybyYF8bH59wqhvhRDyK3PnwBVX3A3spIv4Eyg2rR
lgiGto1M3mF+zaKqdOBR8qk58tA70b0Hc9TOOXgd2eBx34ShRTeTYK111AmghJHUAFax+K5pUE7e
HW8tpigz3MpsS9r08AFyPhTVLmPzPujPsREHtD8c1xqZBVXT2bKTHvbVXcNWfi3VgIPi5jAlxc/q
89prunLC287InqJZ9adjaij8Ugx+AFJwUNxcXhH8vVkxw0knwxbT9YnoNqACMT0VH8QV6VSPgH6Y
VSIfz5roVAxCcqlZhZZVszXUU+urDv/Gwam0cLsua9MCc158IEj80kojsHKphZdetGiDCTddCG9I
1PadpvfVDoRr8w8pcff4vyp7Wc0lMQc4QL9ACChxaKUyegvjSBqJGihOAcZd2HlcilsVOHFf1/1B
xZszZqFBzpnCPrYgVKj7Lf3WaMJR544xLzME7aIb/A7Q9bOSMumkuFT/4LlxT3WbVY//vsrT3XqK
HkXTiQ+srTaiSTw2Uel7zppoiBwFKty9DGhl06K3rnh0Z93yAfn/UkEjs0xaAOxQR+qqMl9aUMq7
WLpua5kYe2nnNvfY4o5PbUEykx/at3iWBymTxzEdlz38mm0Dm/65CI0uZJnOtAV0mcHMJArXLcZR
kQNoLrtcv1FcD9zA2KftnKNqTPqZnw1IECKYl9ALQd2F7KfpFOwHuymbHHdqQyStgHQuSqb8XCO4
QZx7em3xpt56K3mDGmLgLhjtwX5Hx0L2uRDdkxcSjn2EC3vJrT5sszonuTCZz/kCa7fZxk32MzM+
/l9QakMLZgN6Oz9TW1seC14nuQybdqw2I8so3IRxn+u5yhB6cV9NZtz4W2W0uGmoW9B3wIw4XWG2
DYI3xUUkVnSfiT/ALTKRfaGU4j+nInrCvcfUa737KiMM+1AprtC9ZlQtCVLpb7o4Lv2R+WFemZwK
77vGaIMLsmOyTpyIYYZ+fMd+2kSnj9lG7rRrnt9ez6B3h8s71by3hgoD86fxBNNqFOa4BBt98s2Q
rC2EtGbKXTxPrNgUOqzsy/zPey232QtVDcuQc9tnH0lzmNOK1PwpX4EV0E0unnj7uAKrOgbSEeNo
HoqG4wYsa5VZoabe0I/CR/7CukB+H9LIn/nRrQsXqmh0ibroO4au1EW1+ZfoMm9Qv971/Y9h5UuO
ffBU0jVrRdyfn9U3ieo8HSS+HHEcdMtRngyE1j3CkqGRKAoVQR+RS01Yztx9hFQgKQB6NsGSsyJv
mw4jAMV/nNIphVw4nXqqK4ZrgCgYNY7FD3X1+Hc4QFY45g/bO58nDwkSJrXioAC+bGOHBkU2kuKW
FumJn6EAaOyPMg5edk4gIBLD+gs4Yd+tAlyv6HHZ2xuLNOvwdthESbPlzz16eVV0SOyqo18YKuXR
Q1MzkByUU0jY+kPPhZQCsmJYTeYl4B60mhs3yzA3TvaD5Rs5YaVCvZnYuK7mMBdKWanmIHgAXlGC
XGMH2xtHwEHh4gGy+WPFnDi2X5hM+j7i0L/WjBfqw6L9lz8lrSBBy2HhdZmUkiAtMBJb7+yk9nVw
ApWFOSmC/frXJaceAP5qtPqG8t0O7JWr0O/cUg3THo+BB2dsXWXrjmXJQbeCpzZL7MHdQ0ObKrTK
K/eumBJBPddtuCMk6FxS3uoBgZ6qaenZTcKkP5Y0ERbw7QJXpeO/R8u6fF9RcPvDG/Mf5vzGCT8/
imGoWPM4tJPZBgsJKFfzhj25Zo/BPmcWoGbotKGZ0VQXkpAkyFze3w9W7SYWtppuZrpOJLHn7nrR
t8AxwOkiMSznnhFaXojEX1z+HG8G6b1DNg26ug33RuznJ0OgdM/sCwejFxG3GU5aE8F7hMzWbyVW
C8yh3KuhODfyQXdYumrX12ZmwwUV8KDfZi4Kv7BQBWd/EQXY9vd8fH8pgCYSDx7i6wfNBDRVMHXU
jt9ycA8CLpClKrpIb9G/CMFQwK6EUjkTGeOcx0g3b6Gr+I+zjNu3GDJrGOrRYYwXfHUnhBP7PZ/c
lkTeqsxH/OO5nd07XQho1EWuYU660lRHiM4DKHwCHF6fq2gsuDjPgsX3+Xi6UTv6hfLKlqEe6P4U
7YIaxri2tlgd3Y3GCSJBisGZNqM70ETPoCKrPzmycLKTXCKRKfwovM2x1lgQeeuySO3/PrCMDx1r
25tTec7eOHcEcTINyf5ejeHDpVtU5hU/u8PSU8u9Ef6BsJMLQDrZ/J2rP4NUiajZkvj0lE3Y/ikA
6E/p0UhZXvndsfV8yK4aiNLkuhG91mKT92UZnCtVIu5CPQnj2Xx75huJtl4OxeOQCrGjRFzKnNKo
XGPacfMj9Ht/0lAqtT9+VKAvqHHPfrxBbds8OtM698eL5dqrnmDcrJouI/BiN4qMfBIbNIRoKcx3
kYe2TxDAJ/rmmcLUOvV+bSm1d5mtdtTbDFwEogOk0YfOwMMDpKWHyfxXa11N7NJU+9485mbuhWF4
6uBg03PkqkVDXOiQQMT7y7Oy9UtCspzn6oA3VvY3XCQlXnCqBgi7oA/xwWXkj3zWAIngDkntZXJ6
lmRabSsXYZt6pBRXF4qde6tIq2CDOR4jqypeh9L8iC6qfGtT57wHzWXhlSFWl6B7T6S3qlgEjij0
RD2bJr0lUn3Ii33oNBPCH8Hbyu8AI5vQc6CYM4ZkPmndrco7F13va2zGweovJEjBJBSZHVowav3b
Sri9mqOQaNsZzMfaEAY1eVlwnVy1CzcEEqvOuODN/WgRckpMRHJIRVlzxcdBAF+MRpR4ENVyN+NR
skkhKHqw5nfx6neVqy0SpY4TzmXNxEYEtXWcVL9npXMZAeqMnRCsI1pD0Rrn/SJExFCbO/8KlWki
MHUqVQVi5U26MwkfGoG03FD1OsOS/XBEJ86a5eF/71aRPLe1GhTpxld8hsvkHGNTAc21RrwwXaQF
64bBUWEo6Hy9yd8hnwdkYLLxyx92gn0Wt9Nt9RcC5+fxkde6gPLDOqk33iDnP+bh4k1oZAOsPzk0
OlZFgNYy0+5AXcCQN9x1EtGLgkfNQbIqTbRVQzgAhketa9fM4jb1DGdMLPLDhC7YbgvzpFsN9vT0
l0d74tPc5BTR0qbntISRUdI/Y7X5f/0DHddDkI5uFPbkNIIZJtshZZsXL1vt2XQ1R1Cv2zIa72U+
TNl89mJeOhkwzTxC+NqNdCE2D1DwYIsgYFqyPzlbUiLVwv/dfIqEXqY2o9XyItDzIOPSv9oezHR4
T5dwNHiNakCJN+6y8JzEsQsBEMdBkzedLxtX7rDwSzR2nNqgDFCDef8kG2PUP98x/c+uwIE6Fbx3
kHfaQNA+9Xz6SXXinYmvhYu16yyzDu38HIOYimKhMMT8az0lqJTrb+aNfywUwC7qmqodo3jk84jq
0XKE8x+J9QJ9tQ74Qr0pXTCisndsrn3uFnQdx1K1HmjAfTgUH0wnHi9qDElON1nd2CfYuu3XZcy7
xRmw9edenkvKOXVJN3vgMuiVcyfxTXVDaMNTURgrzMwdWtuBN8ZP78d+pAm/oULW8sZ3hTBCq8/Y
o56HBVyBOwFwcDAZ0XQpkhuGfYFjklfZCjfhW9lqjGlUm6k7k8v/IEd9EGEBqILv/1K3J5htB6ma
QT/HY5n/m6xg91PvNCLGklq7MsGalOwJCDKrUKWENpNxy7htPom7CqIGwqAOSS9aazc+CuZbj3cD
VgCDQyk7mQ85n9jN98vci8NsMN5tcMmGYO+T5xtGGv0LaZ3+MVaPN2NcMUJcyp55z7gCEdfjYmgo
mkiRYAc3bxAd87ofQ4BclrH9YBCugkBYoMHL1wp0fnISZzDqT+ro1dn0HQMW7TWjIUA2enuj1gxA
6u0fnnrY+hB/lan6MF5r7lbOUFctntAb1onRlqe23jfptV75A6vhUJ0GEWcgCwbkmKxI8f/o2R1R
lmr4NZRoRrum6BjV6Q//93y7hTUiKWtQXUOg0OBEyhu2+NAwjkB0UK6/PML9foE68F+tiMqYOiVm
DLR6fTVnktX3lmIyjaSENsLCYfAjrw+y4AT9h2KvWcGASARthN7EDn9DwgbMGRj4dcsNMZ0+vDm8
BMSQhUUuPHJlBUEJrcQ54ry28pIkSYe0mrJ4FPEtifm8UiSRldUnM3S3d6Yzqi9pvsrV3S1iTfYC
8Sr4zF4xfmWsZ9KDaTqf+3iwSlpCXz3vO1mZW9pjFfg6/1IJn+YoAjWvCU0cQFpkvv8TofB+HbjS
qLFYJdZdAoaSSSrxWOsEdiMby1JdUKm9FjJX00QfKTfU76rBUTrundE4dfMglyCPVSYyC9DhhUZC
IWDR6ORwUgwiGwuwAXIxobo5DeMgmpCmNdF8+u9u7wkL0e2CglkYv3GN3FVC4H3l+1NAG/t1RnQ7
wRXsifioxp3jW6aSpcJ91aQqoOVo8/RIsMha43YfeWABnx9l4v4UMaCHesjcdN71CXK+mWSag38A
Zkzy0bpF1Ug2kNRJ+Midt6Ll/q2LX+7w3CkwIfp7UXvEodN7dz2FNyf3+YL8ZlTQHqxEOiFkjPV5
OXk6avRqR0figIAzrjtfOoHOzOpZBeDyjaCopSP02UBYMwljkJ4Z4dalDiDR3/ndHd5KiNwCvJF2
eb1iXhjcu6W0YaV0Swtfu8OoDO+jgbdAQ5tEt1MrGGVC8ypwTb8KokXYlN402pK3EdW+Uuv6aMBB
WEtamsvPhDF7I4VmclLMlab27k2tbxaeULU3gJiPFk8X9iu/mMVam5EAz92X5UvbFzwFPR/cEbQd
756PMexbXn2l2s/R+CSiDPG6/vS9s7afieSj6+IDIELpTvtaw2X8RaHr3CSM5EGJ3cNvHRaUx5IZ
ToqxmgoebGyozknfIqpRCKTP8T5UNBtpa4ci1tbw89xYt/Af3rSxN+2yknPHS4GzTQe3kg/yKpX1
ydFJKPXgbe1SlhhBiFEbTUPHo9EP+LH3a6zG8MmOZPduaxUlOxQyf0uyVavOc2WS6ivkXTLRo7hO
i51rGsI4qrwt6gs5JACtZ1+uJjslPpeZxMgzpFgCWZgWCR0QhkqbJVz+0Z7sXDfMHSIVMthPG+73
FgosmoXZ5wNY+BCRWxCg6FhzIAiTPi6ThvpgfyA0xvTXFHcya1Ej+QBXMyt9DBD5X2i3vQBdzEmQ
mZ+5Ub+aKd4ItTqJe7Mi6hE+ALeQIdLhWPDfZGTLw4T6+EQMNZkPLd2i4gkMTFuqH4tQVvYfhXa1
zPeJFk2V7964PztZ0p0nERaRBn6uTbPv656/2gSMTeoY0WJjEiaQbxJLnX4D0gXywDfZoxKdAQio
+zaMoPlXvNHyjSBK/+WfDz2V+potTyFgfoqR5iTz0sK9TsAKnfNn4JZP19MWIv9QfgSZAgJB4aWN
sgTVpCaD1aM71hp+kI56mB4mhFy5LhTE81fCHJJ3DNHOpP3cuQdHqDBgx/MEGDEQ/na+W3uoaICX
WpJXulDg/oL/dti9pwKoWH7vlH4sX7TZTovutUw3cwCwRngnS2rGdwlj+8uFjnGL1uf/IvvGRMy8
HYp73Ea99TefTbTsOhQI4e62WWWUvPjra6u36o6d3DIMB1C6NNsIf6+h9GwdspUiBm/qPnOzd8i5
4rGib3Z8sOZrg7zSEreez7X5x2sBUpC5GDEb1gzR/+Leh+a6cMV29G+WNcMkzD91Bg/a5oHhVfB5
1yezNpLZuM/Lf7GYTSwpHmdFf0shiOE2gsBkPrJrHKabc8Ew4CI9JkmOl0jjYRJJ+Bprz2ypMIO+
fhYvx0a5LGvqhep5qBtuZWIilodnyGW/808xgTlgpYLKrosAaUNJe72ghO2sXAe7qptdbEEoaxD+
06+uBxcsIvRHXmqqEUnz8i+0gFxtQUHcZIzYAEWQnVGZpFSu8i7R3+GptsdAP/9h7nNMVx3NfV1e
zcFFOdOTRImazoW86mMZ0ebUxCOeCYu7uU8aO69AkVIFiyY2JGtG4rVUouZZyz1mjkfifPYN2ExH
q4tS4qXBNe8lfM6EQ0VwK+9Uxcl0QakZnUngW/pM1YLFQ/L1vfSrHYOSpFN0NUVPdheQalSF9S4j
8eN1Hlkj1t1PnNtIgdS9tNsAZzh/DG+s1ub5JfVmF1NKYigCzTx3WKlZAkUCJ276JAHR5DY9QN39
876xigEQh9yt1kqCQVaWLcJn9U4TAyWQNHEWqPPP4F3neOvGlbvt70GbScRo3owXLnQ8cJZ2PbWj
BHWxx9k5c1x00O23q9yO/zfLKG5a21d5x8EKyPHZAtIMK609kxMKrGp5+leQj0RHph6aKkmQGhv4
tTxhpTYq5xRxPWFnAIJU1GVhvcptv95MW+y1a4QESZ6zSBj/WOJHp3eRFm/XCgNZSTQh6WMk7h+3
E6ulo2hBGFs3dicUqdd4r6LaVjSCElTV3bf7dcCIQjydRcHCRfLWDg4/MdgUS47x/Vq5oW0GkVPd
aQniHCflp4Em4XWk0lwrG2jKDpOjR4EjWVPnYrNnxMcbugGkzmN8jh+s9yCOwNHHQQYhNy4tBPqX
R/JRogAmizcTuOuD4SUk8rU0jLLPqkNH6GRr6Dtn7D1PN1HGPcj7RNGi1uRGBz12r70NNikfoO2H
C2d5bu3hJ6m6anP9It5fuYbH6u+oFfLeUpjAiAewnS5N7CmtraIBv9nckPoIk828pK1RvrTYc2xK
ezvn5fDyUvaI90VsguobrtsEe1YFBUk2EZkGM7aPmaa893VLAzeMIehaxvm+CxbSTfmDNwVYOYPc
jqr8L82Ewvvdeu53dn7T6b1a3ulrqfyxy3sCchaiAMdUIK/QybLfZGgZZasZgCMazZ+LD9sz1b5j
pMZPQhN+NnJwOQsYHZLeRUOPodHJMUs6RqBHRHnN1elEkgLMQq8atghm8nc9vA5Wr7uuK/gTdwKM
3/QsxpV9tUIcP1AKyCtG9k/HOlSeMAQxjF2toJ8ORAD2laTfhM4/G5bcCL+dS94Xche1Js5ezR+4
LpVtzUUXHdx/ygoiT1irCcigol2GLd7+WVP7CI799nlvKlvZ6gTBBGRbzg9LCffjafIqGPFq2EvY
OwGrNancr/644jc8mgLgm0j9c4dKcxK70LUyAVCnmH/v6kBjk0ijJc99LsBXRHktgJFdpytJyzuM
hLW4nPc1UjHSY6X1+V5qs1ANLkHJYA9eAmxCHYHkVEFNqSr0/cK7j4K0yrR1jqFVSPCewVffz60P
ufATuDZxTAztPt0Jv6JFpJ2TRMT6PViHYpPsfh0J4AhuTFBhUMwM3g+U4ek7w2QA2vmbtlezns7L
6LMcNydXDN4cr4TskmWlNBpRrfI6q7nPe7+xEcec9SSykfFCMc2IgoayGgnZdcaBlAeO6gmYVvCm
ZhQtRr1l8tJSTEDkG2soqr5V8Zl5iPpkSNNft/8XYIogCrbTsEmCb3dCKxdBQSn6TpkezjrhPn7C
eIwRO+CY9qrSBx8iGVYa627dLywxYiyPhqXVdpmVaeGSwniZKgoZSaRxih4K5j6TVZzI6Jp79ZBQ
6yMDs4JOVGuqwUiGPGLWqwhySe0mCzqJSnWX00UDqTDO1h3lKxQdK8Z17ypum68bTvyEc+BtrdSR
qWjD5uaGdNMONnh6USjhlsFKWKdDRyY7rDZkzIVVEIXrFn4S+4iTbwUJZVJSIz4E8GynNYgUjfRZ
ssFfjj/UsjmkSZwc8vNcg6KjmgB3PBnG2qNn8/vnLW2KF6+GmpC0WxqPkECbusWFn3N5BLoqYpwK
vZx3Z3q9La3MVIH5oQgZdEvkxfuuZ4xtbNbOp0rp0eKlnocLvO6G/bLyvqoH+7v6XmlOiFRtGe7b
SXh/bEOlDL2zcja2beMpcxLIrjXg0rnQhfQipkT+f0er3T2OZC/fTfdLTrc+KgD99jTCtTAytloK
GzNFihgJZbD4WH/U24RwzVQAFgZ3SYSnfQ1+5JfYkl2PwVmrJE/smrULG28aymtxKDi0XtVX4san
8+CAzX2hnd8mp1N3ruwWywmZz6PQgERYFeupE4gaG+JjsKnuzMrlZJ4TUN7CKY1+yv9FjiZny+LE
Vdz69///3XZ6FRO3CdWUbOMkJAVkQSBWYp/hH8/GFLZDKKbzCPMNObfpYX5Hz8XawZAUMPqfvhh7
9BhhLuaowy4k1CJFrv7jBMhVhxypBx/cFCBXfzZaUJzseUUIuh2mEI9gf9+1pyJEaCTydMbKD4e6
Xup0bSTD/7dVCGQD9QQ4sZCkkJLoi/+Gzvg2MvQZ4ETm39SD3GCqE492Ic01ywvKLglTSh2Zfi8+
21Bf5oqkQ6O1vSpTyMaRi58C26Dy5q13Kon/ZihtYbQOxLeOgjWYhLgcumzJlTE/hLJ5ktXLl8BJ
LD0/yU4yZQruuSVIZ2VxdU9yJBvPkpFzkkMbZv5cbkKvtTkZqJJhm4LtSFTf98ogUfBZtYkci55O
c8VtGFvXutIFJQN+rhVqYMySveqrhKgwHf+5LrPbOVbmW1WRapVRH8YQ3Bk23ErvGxnqCDDssdu8
06/zftydzC1vT9xXQKg1VLv0sUIYZ7AuDmnX2zBFV7FJF74BByZXqeM3AoAe/q34ysXXfk/y+ZTN
SEegiYpRo3Xw/ozlqwrVYcy6c1HdmRSprn2mxdliRcX2ZtwnpHPAke1iWh5FhaP7pr/SJTXw/VGD
un4IXzkCjV8+sKkRvvYL5s7u+FJLq+wORl9bRYZHzz/LBQZncG4UEYXfiCx1Z1D6dILG39SmnrRm
keefoKaSkcQ30YznxSM+P5UTP11ps99C2Pi3ze9OlLnVYaQ39xE2BNUGYVlPsXrqay3pgActgls6
A4kkKgkWMUBs02+7egJs/Me9wJOU/JJ4DIhkyW9klU8g96aExLSV7lTR3d2LZoNyLVHHb1tGZO4u
e5pl1HZrr9BfPWu6CXdY2l90+rQrTWeH7sVXeZH/IXIXTChxN1SzTujHw7IDdzaIjOY1SmoYSKiC
ljj92Mn2+n+BFktUpEU689Axi64QYxWofjHSyT8FGcjxMFU/wM7mHOVgKaN1sKj1fcJ1/ikrpgNl
db9DzrXXFfelbVBKMbtx00cqZqAfeL5ABtJCg8v5h7C8/31iqcBPGmW0q4+NOxEsh94L10T6NOkM
HOZp2isaJgtGu1ipFrOqWrguO4zU7YVE9uDk8KzIflbvPBtcZ7tVVGnlUFKTEEgZUHgNWvLVptN5
RxFDmSNoiAMTrwmMWg6lc9AzrH87eHSoj+dQ1lqMmzV6Iuk8Zv/b1A9gFcjxDjs0KmLc9dY+pXpn
Jjb4zMApsHkP1CcoIeKVPAU4Fs7D9i9IIRjXJDkaljMfTCcfEne97UP5AUqIft7xDvDCJovrbh79
EqCtiEh8R210AOLGyIVRPkteBSgY4ItrUoVbJ93zuAyIQdZprlZWue+HcJxTJwCmubXVqiLNxzir
7spROZxifod1tvdas2fKkJs1vaWaCdeIgXsVWok4W9UrS+2GXPHHpea4K20T3ut03kDg4Djlz21b
LkrFAxYqdpSskgBzrtGCZ2/409dOxDkkt7FSksEJ5e4M8ECP2zgUFqPhq+6qBcVGtqBvH6urQae1
6ESx/wTHSNODzxrYrMEsXHKu6wUxZWUKWy/kE0zK85QfIYDkGZCu+Q99L1brfKyZc9fveLHll2QH
8+SnA+VjNgm9E06H7O+phafC3XxkJV3JAkwwuETm5AFarvQX9zNFdtZp141AM/ZXJG4UzTBa6/Hh
cYeGAN/9JbP4PnAsotERdGH3elgz7p2wrF73mNqiuhKbRrKuYkWQaf4cKFVaB6KNrloVieJVkcTw
GaLDJWLKZ5bwP/2dNsi6JbKAHkAU3wn+lMn68CBgt0wzHYfk0DA8TUTdz2o1Kz16PJOY1mtnQT6g
mRHFMpcXonU1lt96hKOisbjIcWXIkbRBrWLnHaYmp9qOqrhH7KT5asEIrXj9OxLkAgCpTo/IQpCE
qbGItQFZHpgr3/GrA6aqFXZS+rhjysDomn54+31+UbBg2YgZRf8TLHYQBRtdSmDJCDMHcnBpGLqA
N4uh27ivOi0RnoMXbnCWgNSxdORcbbeTVBWK2TLfIvQ+3AIK81QP4NDhEsX/waOPaEii1WBKY75K
KBWiHgrEh56abYvDecBWf6FW2dWVInCG5HYGQEhtRyYOac22KQvLSra5xJuo+GgbrcZp57fNr03v
SUbY8NzAmnIWxyagMX0fr8VVtap2gmJstiewGVnsyxeHj9/sVXysLi/Qru7pk724ZWGLAKUZ7XGJ
w7+vShgOHlBsi1Y319+lBLFwgfFCfsrqJx6P7pAc5AKqt0LhrYCDFwf0VtxbYOIoGQR207jv3zUe
wZuWGpWgYMQ7mudmGjacEylTb4SsKMNR+ro8Ge5QmlEJh7iz9Z/fGYshIytgQwI/s7k1aQdWjHQN
3B/+RqHCQbcWIZrIotPsiBEUI/n5nNKLp35awewMNoLgR+/sdkKTY0ZB06WpSxji1yqImBq1MLRp
orDvCM4xoo9++Id5xSgdT+HQ0b2DS0YlkNWHH5/LI3oU2nO5i+WBUqwp/LhfCPBuU/xEEeQqmWuQ
CNvAhZ5sYiOxDHqhKa5Xgrgjfq+aO/0UZvwD9DPqGxK6MG8f/b/Oo3hl+WH2Z0b9JtoEjfv2PgxB
b6BDWozMh5h83X5Gh2cyygZqmGGmTiBWw2XO5nqzH5yFFwCLDvbWaTJ+EBcmTCr97Coxe0+l0uE0
V4aZkuHoZikM5hrKKR02g6mQsbLEO2VEMmhJnwYWU3RVF1dJDCzTYja+HT/W12hKszHjpczCnMSG
1m+B6D2XJNuMG772jx4Gd93uuDvg+yE2to6qCx1AZqZ3Rmdhbe3XIL2A5YoD2rUozORxwCPh+v5O
/sdb+NGaw1s6H/+LRezZ03VA0AANG2CcUbgLKCZUFVt8GQybhQCcR5KMtfRNcB6oX6X/ZK8tbXz9
QxkMGBQvgRQQyfFfWzE9mfVy/IkmSx2tRxykeD46suHrVDgyCoO7FDDyfi/NZ/Y+AarBDPdVUOIy
xCG+177SRY0t1bDB5ueShqodt5sgs2W4Yg8vdHV/vY5x4O6r+F1YKXGklj4Sub20PxOrXmamuWia
GsW94ye7B2hoSRSNWSXQ58tENM+fOWOfG1lDs/t5UIfMiWeKkEfRiX5Url8p0DmDL8jX98iqXVfL
FhuV/3hmlw09vZaYxsA31nundQ18woa4Mcxk7S8NTO5v6YSufiERU/JMsQBQzKhUR6hMpSwR6N/T
wFIgTRYXfXKJlJZO2/5teRUk6tKc3WzJtD6+YCl2cYdfZoujNaPqXFHxq8sogKHzxKNAJhbeEyIu
RTqS+XdpTLLu/hOYe5Ujv/OUP8vM0a5cmtVW90QM8Na4JvQPck1wFD+6yvYaQHby05RmwYakCMtm
KeiEXCy6/TBiTB9voynMJsEGApPKN8tdPw+evn11rgi6qKFVCOQCbguqh9dmVjo1vva78+og2vhi
Nxhnq8bA6dAsYgNDfLmg8EX8xuIIdJIjKw3rv7/WtscuHykQ93aGrWUd/zvoeGQv6BFhtH+kjJiv
4W+25bqDpROJ9Eumf4PHUy6sN0GwdvzS70VTUbzlT3i08dMfo8e5vLxmBD3D59Tw7//PCJCJIjlr
td/ikjenjC45hoX62C2TLm/EiMQhSO9jtZisyvtw0be1BQLwXcd3uPhhx+wnkrJ/wgY0GAKVcJ2v
YvAxfIu22Tk9HTEYHOhBQkIGkNmMXMhcwCZH1V0Ms8VKVGH/xlSVLVV8AOvzyhX7rmSh7vMrWNAk
OyqDwc6A1mXitMnk86Hb9kh16TyNDbGtKcYIIo4JPgxkcjpw99CPa/EUNRQd2dtjch8RXk3hmgcU
A4cI6izvSDHlsdhzWfRMgpFLwO0RrpTiP3MlUSCf5fgoPn2Xxcmnrl8V0JvyZXJtKsttC+JWhKxP
jfRZzfykftSzGRVghVmz5y2FwMRGivWKAqQ/Cu6DDgPC/VvMe8N6bfyv9O9/Hzt12r0DZu7r1Xgk
9dtmnfapMM+XgrYBuejFvVn4ov3SFXe+IzIxLdTRpY5tiHfcOkJzkfqYTfOIyAp2j9iwSmZc5aLb
LJq2HP7S51r9vVLINC3DZyMXJQrdTd6h8pFNg+dieJxTvQ3Kdn6iWGFr3Y4jkqbossIdJ/QXU4xD
bZWClhuIhH/cIieXh+aEhnbnLstWj53ZhmPPzCbDHcu7aIFNgfpABsBMgPdarhj+Ond2Jnmmc2Ta
ThZV68SixksFajDvyYusP+dB2+SdMEdy4AGkB0tNSS4yPnfVOl9X5mPrW3N3jvS11flnGNtumbKt
6iBkNxewooKLWw1jNqJoWmmVb7DB1JxOQw+epibRWRCFhW/O9+X5+oJVE3L8UV91G1YD3GFPKg1g
FclNq6qQ8xmPsgOVcNAbPJStPz2IXLBtR9FHtaVjtjIDnYSWdX/+YD7NJdkedgEvtCbDh8nhzDos
tPKQ5H/aN9rK3k5Ok4K7DKY8miSTvpcWtLAycX/qtrNvq9sCUrqcfY4PYp1YjQJU5x8N3nJI9B0q
qscxDI5iauYc6JxB3jKtuAcgfQx009EfrWLHCYOFxQp2YhKXiJ0BQ6S8yasin5Wt59ceHNbMPhDw
B6TJkHM2u8REeBWvBJAv4R+qWc6SNpAn4rZnMxvP4HKHxv1gLXQltutbkwGwqjqpaUNLyusk3SM4
RUd3+ak00vk/wdsKr69grLC7FT+fUvhFpmRsiXkKbBiSw9hCJi6W5qpiVEbA/Txqc1F+8pF7GGWh
NxXjm6pS2W9qBWilwn9TGxvDKVEb3qoFPOohIbmdtyldYzr9n0E6c5bvyxcNHKIhsnqL3QZWy8I8
u9SpWNnn32RTp3jKMI5cgAdDWu8VNB+5n0NnRnlS6Y4w7oUCRp+MBkBdmkK6VkhrATwulvDW9Z5N
/FE62MN7ncvbAs44jRq/LEjvDeWP+5TGIR1ALHcZG8Qqx4Xm1600OiXC5NjtcP8XF9uVBB0jhkhq
agoC+oVjznQg4SpVa3+/1TJrQ1a416veKH2FYG9Mic52cr3Q47+TbhIYdrJlmRdjoJUlvhC75Nz4
2CCIeW9KP21r7Bisj6AkYS5Q8ehjXI4mbsY4AkngFrj44H3u5AuJGGiDNklPmgd4cR9LpgvrK4oW
XqcUhwwr/8qLDbNhmZ/NX8dOjtlnu1H764y00FydcJC6xfr89/7R9rULICX1vgVfBYMo1KqIeqTa
J71l3QPp/bLFgWz9SMONnSeCyGJc0oULqfrUsg5f44uoWCxcfBCRR4JQqiBuQ92wSUMbdGpKiccJ
UYDgMPJs42gNE8fLdUDlMNmH8Hb99ZgOkFjv4bYe0ijR8igG6mj4zxKuT4eu1eb+ieto+kNxQrWt
cNNuKGx1i4n/sLf/vw18dGJ9YtI3bchPYhj0ozgMBO99LiFoCAvWWbiJa4h3okRP2ufNHZD2lhju
9PzYZroNV2HogJz+XnxhfycsTrXSEgjl+vyvu5z72ejuvKsnZznoFUIB6giy1C0i6EZ8TCzg/IEy
bFXWQe3nk89Plu1rYZXO8uRg+GG+fRF34NHDFfg2EJW3ruNooKwZI/pj919tiG168FZSS9/WChYd
QHqsMOiStCSXDoCPm9HFf33pBNg7fz3G/254yG1pKZ+XNh38MQPLnWkGtIMhkQMxulJJODogUZgH
hM5uw6CV41N5FfcsIldsTGZp+NVOWbP4xs3fwYNQ+xQ1tiy8ErFF2aF108IctNLSJT3qtMXf+iF7
W4hzIyrL8d2NJNGM5WkXqKD2MvpyNfUVTDo1OB3jWoNFzSXby7e/eRrhfWPAqsPiaDWjt0Dc5LPc
n2GcqX++PoFph82YIBzcUfMxwAGF58HCJHvLQqypz+ddGKx1dT3LRBIlWv7vIx1XPWISrE+oIPaq
h51AGyhKnB1rPYxhApit43aF02EY0cbR1D3TvJGUCpBiquZ+QM0GmxBodJdckw9qPrpPTw6tYq+P
XS8Uf2aO7iRcKcFSfHv4eZmZ9c0KEEViT4ZZZNGhmNXPaYtknBbYKKJLX7k9DLvPPul0qUWOEPmN
TqbJI4NXAYdZ2JfSjayc/1qk4M706Q/kHmS+BZx/bIFTB3XmCUfIwqU46g7PIa4T/93VYP2SISAw
gwMIePBSZGDQ4Rv68L+/+DYIGRQa0JQGHJSBD2fVSLvDPPYxk1PpIrfalaugQ93BOUTxVflbp8gT
SlfGgBZjXoJ7i4cZd/Osiihu7gog5oncLBoLHszKHA3RNJznatCfFLPP8407EjguF4PIaKJ+co4D
vR7AETHfSVty8JsRdhW1tw0bxANhZK8Z4LviirFMiV5RymP/oD21SIwWxCK8ZVejx+KGOrA9H635
k9m+7alWb5b/irPGYkDkErMvz2GDpAWhxO1lKmGZVZ/RC8HApij2NUZVkMNPi13arismBLPXwM/N
e9lRnJOMwp8+M0vdfOxol94PUL5l2yOPnR/Pp9QEsym40sr1ehbXO96nf3JaHkSYLs9/A8W2HMA4
h65UUJaoRH1HrfWoHjFo+B3g3AHA50Ivhm6MlgNqZFQclRbmghtwsA2mIxDr7dh2T751ok/l09dU
K44tRq+XdLtUj81VTbyg+Yo3bN/91Dbo5rvOHWd9GVqKtu86wCb7EK6kBUaUdxhrLcV05O7DHUVR
+CdJTDdS7X1E8Kl8wfprCSzEKP8da6wPKLnBgNz4IHuqoZY5BakOAxe48KO7C3Yqfr9tbDcKsEe9
n3G7kQ/B4J4hqtje5/jDrjsN3nBZP1GpbWkTRdxTW5qypTOpX0spAMfUrXsqO3joR8MCSwQRb/SS
EJjPixBD0T3dSTEzFUU3mM4M//X3/jtm1+NXowFPv+VcPqTf3VudzBL4WoqQReAZfM9Nq8sdSgkp
1TWL/etjJO05Y1UjL3s/ISFSv1KePftkPWpnIZjIBfvG2A9/25ruPfCXb0YnIkcylI0OUJcq/93t
65OBjurEbXMzPWSJbxQpPP4ORTXdlx2J1stoGv0gGDo9zSJmK78Kk/yt0ULYZs0N8ROK+BVSymvK
8IRB1R27YCL3jxK9D08xQB2q8/hLTLSYsG0lcpshF83aRbUajm00SCP+PTn/GO/btaav64cUMzMP
HF/xyLCrMVUh4+ex1H7ectVPe1ri3QBWftc2kTc08VzgzYlfzrP0oBids8T2oFLkBQaY4sy17gFK
bsaw9oB2E+lB96ngSbkyIvJdiJP4HgXSWw5UyPick+PGsfPSz5n9MTIeodD0k2z0vZp7setOucwf
capJs+nHF6aFvC+/Dc0x3F6utqaNi8gMnWQScR4gexYFddK87JHS3W0gO48MDVSU5GWL2FAx7cDz
zrwL4Y/ijeYBt1DrAXNd6bRp6Bgd+0i27Z3tsf3B/WPGBV6KFNaafRfg7t7JHG/7KjhppzGkG1Pn
omok0wkGarvYdG/aOZMJLQ4+lUTB93zhT1uEFkvStNUGD41i3HNviBXT+q0wEhmEVAtKk+dT1dFQ
Eunsjzsg4ZJ9cCDEQsGcUaL4AkBLqjPvGXo0A1U567xAX5Fl99oakqZkLn7h4No4Hykj5DCmsx6Q
IDUb32WwjjzRoZ7tTL8IMSkLnZ8T20GjejqgKsGI2HLxDuDg/wWESK2VdM08s+QmPCQqt2U4IMy1
dLVN3uZV7I8tMTsS1ChMK2xisPqquZVxkKfKcueZ8zHoqwjl4SiUpcaH1wGYLLB0Pie6fcrCvZDV
MxJrvTR8VsNNtRWX5DDliEqH4SxKa7hDCHnLDd+PfMlklkg2E6HI8MBjjt80FBA0PvNoEPzlU+lG
r6jyu0RUqxurXrDwmuw8zDJw4EJdwQTbVcxadCRrdIU3WaQCKXQk4+8kX8fAjwRdse7vZ9qd3EH6
GgcC4VpeGwcm9F9U1iBF4gFDLAo0df+JBnVAhdukg9vTmUfd7v4Rxr1Cr7miM5RIWYbHLYsxuQdW
25IokrhRqP+rsbeH4FjHPUeciLYK9VIjmMYShSQHFKNPs5NvToNIolJD5yOG5JlH9SO2k7TeV6N7
36aoC2xSE4h1JWxVcwKPY04/SuH6DDsitwQrP3dABxZUg7LxjPHaP3x6TMnp3dP60Fls22o138wb
aIM+eONpDlDsd4QYYZN6r0ggTWWBQDGG39uRX1FzYL7k5akhYRWumwNZkQSXBqsm11BFGBVgq3fA
CRMuORsx2aKMLOwxpqC55hcl7n5aiDZ9RtYOtmhSGw7ktmwM+r8EJ4vEpKlz947DgACpFG7fwbcO
/YAHuG83927QfLiy7Ox+zS7S/cWXAKGPCxTi2sQWPA+5awl8fG00atVTTgUwIItMRet7zFNprSfo
Zk4TTKAZzd9uzNo0/OmZeMppfEd+UUDKh+9rKof+eUxPcZnerBPMixw3PDbk7KJcKAu5aGBsXVov
AOLLEPMqdu3cUS54FnGrQ3/cNwfVdBZxsU3AHEJEjkWpcobzaSMfynVaas6FfzvIgTMYPlDLvn3O
thJT9q0r2V2jN9/NF6gjOyw/INPbysGtw5OMMLrlI1/l2BJ3rAw6KePpoee/7mBR06uQyJC0194+
U+Bjp6dvtSqvuSTIw7EtZUoZ3NpjGz+67mMzfhBl8iIbSu8nnNyvxB/BhwLVDeUSEGoZ3FDgdnhh
hvRQNjRjT2NWpwTtdYwzFt0qVexKFozS02dIfAaqI4/kA7ubFgRViLVMZJy1FiPVkk10916nGgV3
tz544806f72N4EyRPYNR0DUAykMYfxbxBArMRxNvmtaRD02msNTRCqqXwS3FlaDgw5V+KkxZuTpK
pSFhcZVEncrNoKAstTtBGjPWLYTxAgZ5SH3q6vz7/1J9EEN++ysO5WhOx7mtD98pjfxTa0UyraZ1
7lJQZz7twmDOZuNNKmY1zGYRqbZ0Qxt5hy0b7Q5bB1rnYh3rge3vvlxOMwRZ6p2gKTsugxG9ER7Z
FzW7ClRiQXygPTL0fyfBV/1nNw4LyZE5HbE2VWUL0wJ9VG4PIUzSJFGFqy5G2dLjv+RJx38XBqql
sCo+s4Q16LfNvCjPYvfyqePvc1g1PpLpQr5sUESUFVrmgRuMekFCqJmOSLFavv91vnmApdkW+P6Z
FgmB9Bg+Rs9GfQzBaNr14ILXqRQUOGS0m0/sXGZ3+myiQHryGWwr1X7ZAr/Zo0VdS/boRaGLYr/m
1vjhrJ1hbguOn7nA+ZFzscjWQbwFtVoKUR1aDOQxax7vhKeDUeyluGm099I30hwAJn2snDScxt+e
9Y7iOIW7gs11AQAeg8AYJfLTBRYBsTPOqrnuEeCyYnwS3KN9pet3+XmejeiReTBCy4UbFiRpCeiL
gq3BV4Y3EhGDG8MUiqEePhplX9oFic8mzKq1zrHeHCwh9KX86xlvDjnP9KT6mGDjpus4aTZV2vba
I934r9aVP0kVCZftY5h16MHafWOmThNDhTJLRzcCsyXIpY/MMaStsffjLa49lYbsKl2H8jgXX/Mu
RuGUG5yTJ9cl/u6j/dQ/00B95XySXdwtauy8uNNz0xbPQbNzeioy+etK/qd5LIJzmNJ4yilobFS8
qRuWQxTeNUQgBB4zS4ahYSKXWhONSQtmug/6gJS2jj+HKnJmWAlstmrAJmmyHJTpiubPIUFWi/se
qm2a7VT0ooamm9UQ0//ti/z15izpju7FspexKGEZG5aEy/adCtFnSkCCV+Pwlw0FSTW5A0aFdlY/
trVU0Pf1y75QdMNPKMYO+T8K4HzxWcGwAb7Jrcf8HBJ2e0YvtBG3qFinVq/JB8WLWujlSgDE65Ud
+7bcs0AYf4+TVM/8whLnqz82KN9nK3JCENaF6GaFufjb7VkBNeQapiPr0gakMsbZUPvHCKVSf/KZ
U2iC6pH0Ol30VdlyIVI6PQ8mjRow8hGWVNFHfpusZRmViBoP8NjxNC076snVOZqNe0vO4/BMkUBk
5n/mEz98EQ5+tLr8Z/KucIZybdB5sjPf4DIQbCavpPw+km9Km4uH3WG+/EJBYb2koaWJGN/c3dA0
8Sdr77EDXtT1I8qSGd3l5uvc60PV2AmllaksDP0CnPO4+An2sIJDIwIKUK8mn9azJOvstMJZDZFP
z1Ysgpag55WHLfjcO+eLwnc7PNtfwWSj1hrB0f+U4NS5BP7/M87T7W87apD25ok0jWjD350ZGkLV
jMevU8hWeqFcExG5Tfo71VG1uMznQb33T5zk8EJ0hvohpPSMJ6QM0r3shRrAxZ7dS4nKejXL/VSN
OLADCPa+xm1iS2few6CMntnCPYe3NAojyamoVwyO/edgdVkj+6wFDAdcGs7zXAZ2l3Ae66IuyUeM
JzCn82FPdg5GgafrrwjIkgtK9VXEAlimW1QlyXuXcWUbpJw0pl0/qY5HvhhNL04YqWLysG9+zpun
Qovr2wsdk7Vcp6zrrA7V4WcxJVvhSqKH9SgyZtWdXpU4g6JmjDREdO6ONqQdJEyghw8oxzPTpqZ+
+QVEU+9w6/7MSnZGU1gU3CJfwEMhS7l5PG8G3brrX7SwqpKkP3tzCIYbmhJIhxjf00X8FWTqDXhc
dMb5QXf1WnIi2vAMsjVPq9rmoc1hRTBmvnJym9qXHWsq40i3j2CL+Jvpouf8PS76YchMMHLkKTQi
PHg5traVo3dE9PtWR9IPzjFuS4/ISkPot78nT2kaGcVlc9x7qcayD8lGlMvZWSjSTTt+lstRaKx0
RWuQStqL5k+/93ndvJgEULnM7FfaLD52kFzQld8GaiQ5Su1gC3LIJCv3JHNE1xMhxsNYcPSUMknx
zxrRh/3c/Krvst9Fk/cyMnnhWqVia4C7xpI76q/lUcTjUUEdGCh/vkMjTlsGYr5xHALk805pC6uq
7EGgrpDT20hPIBP70x4b7IlwZ+Kt+nYXlIc2mGK7KJbKnoMxbSaNSqZCMpSu0b2F0uB6+ZUBEh8b
fwFA0QEmcxEuG55UNwzN4/ALRgFi2lgjsu1jSjbw2Oc3SK00QPpI+mi6j60DuEwUHZnVcLxqwtBN
fJmCsOoMJgtaVglfCtP92nHpd2GFHHPVpMLk0yPBX4UBcWdhAHm1l8u33SCecdqXKZ3S/1ol1xcd
BdR7inFdCUzGyKUY6lm3fdvCA7kgAngEbHEtT8+9/R8rnkJbV/xl4OzSNfUKEZ9fdVC4EA3a+Xkn
tt1HGTpPnou5UI4w8sq9t3PI0g63GtH/zI7k6qyL74M1KoAdDErO+56If5rnQ3/xkkDzCcmCKz6f
5FUCqQARFsAHOn0ll8w2O4Tf2HOGOzg3yDdwXF8n/O7kkaJKloAL7Cc9j3oZgW3yhk+HO8SiaJQQ
/PujTmaPAZhqQs7nHe0YkqYoN+KO4SCFsW2pHyX+zMWpC4uHOQNa0t2kMNBGzp4K0W1zYDK6nwoy
GV+qYL6ZOe6B75vU461mnIBSHNAvmjBybAQ+1JSapdMumr5OSKLgX3pQy33gM2WR3qrC7SxO+zPn
O0uzcZY1919dqD/n3Zhz/40FTO5Pp1lJZDvt7gZbcWJ2/o25RZmYfczUJh46GdtI9NJiJJGMz/9k
H88v5zxDoX28uPUGAbLAaqAnTHITfO5qdsodRxPD1Q3DW63+FBFZkJJ/VCb2m6wVtP5/tDzd7tLx
tpCalRDmB59Uy7SN9msAAsn7nlCAeLovRHFnpJhvYwrxmLpLiQQjQJnu3od+zHjI7Lc1a6AbzGQX
9DS2nDI3Si3rcJYcfg5YnEUClXWu7KvLKE6RDUJ6rQFQKIQbR1krEEJrX2hr6kenE3ibTY486VVf
pkdyLwuX+1HxPelg1P/RROjOC8jd4Zbi98fGdg5hBoN/gQFwnxC7gBNbvFYayaOFidKpB+FMLPpe
UtlDU0p/PZXhts0Le8fibqCSu76Qb5JIp889I+mbU3Go+9W8zjRUjauiMpwGg9/2gqsMzqEsUNv9
Q+r19ohiNW6Dyf3hIsXRQv7J0W47BqVLXAx0bV5AXkZX6LJ1t27Y26xiRX7gRFc5CGe3ch1vy+6S
I3The/70jjnBCo/WPNkU4+mICqRTVRgmC0Eqb6+84Pv7ClS1c59FKiy6EH8J+PvtcrtofhIgV/od
5bSyuB17MR/sWX4so4Kw47PqqbZjq3EKMX59LytlwF5cHsS9p/QcxGP6vQiEXTxKqGZGFWScyNPY
9SxUdE5/Wq6stFlNC6iHKTl1PyndAW0gUyPgt3reHgrht+UIrSt9f2WbukBab36su0PhzrAhcuZQ
uEqUw23rr8Nlo/l2XKsMTsyWoVSCr+el+Pze4sBmCsNE6dKRQFxV4ON129CbX2Ihzt2JbWIGUSam
h5ElKRN8XEN7Y/v2O6B0YwyQ8z5Q+m/+10/rKyP7VXcgOzy+EGnAQ8zGkKPuQnrxoV11UGpPkF7l
w8VdtLJdmHVpKfwb0qY2q0MhpoXN3hdvqy/ubgIFpGKhZOc5sj3BghgeIvqIfpgd5IQ8f0dDU68l
MxNdXbyYvCzFLmiaV+tZ8L+mKY9/sMPGF2kBYBN3Z5WeJX3pngKf8sOpyrjcCUxjW7KqBOgqmQAm
zjLAe43knq5vnXTWGgN2xP8A6SxPnVYENuKyH46ncVqJLnSSRxDAq7aoGbsyT5gf81KjRSi1YTiN
fITZtFZ6DaCaVtfb8UNtEHSfNxAlkuvcgxWQOWf3jNU1WTeazNzWpX7jVKi5NBOw32diNL4W2zc1
iVVjNAeml9AQR7V7pMLqsatC8WbxBsd3bO3RoS1X161Avk1f0tfIbYV+zihTPQ5I+dC+P7cursYz
XXB8OH+wngYGKWs5/uigFHG6GKPonkXSf2O/khATL4QfcysLmG3KyXlPm8mG1CnM1oqa80fPwEk4
8Fsw588SdOsHXQrZpRpb2YBzUrn1gsJysmVus8AgJ7M0gf12p6GFrHBh+pPyTMNqhQ6eA/XNNMS8
1/sHbh552vIKuUiG9IID4QFFU5G2IUQvrILQo162tkfDVEk5wpvagidOFgDatv6Yc5ztry20fNY2
4XHQNEBRvc2CFp7SkFyaReLZBTgazAjS38TUf5wjMCUtGk/0qyrKC9t58rc5EWZ90YWFENq+HCVq
xlcKtSIX7X5xgsUMurPwntMBQltGGpYUsZZodt9GkeuMA19d+0eTjKb8HXoN1MR9n8JihJv4KDdp
oCzaoFV6VZNrfbqeCtPJ69rbTCOVAYiRtrPL6O9sEiAkbT2Pw34B3PtdDDJVhYYB7mIrAaIPFXAm
O48hra6eXW1dnuLgIO42NQ16bMtR2qqxzKlRO7X+Bt/dqXisyRC+CTyKdbhl0T3IC56RxoRS/GFT
vjFF2kS3J6d17kX5fMbTBJJbLp8HxhYbhL+uZljYUcUvtn2VY+APMQCPOJ6q61E3HJrjmBONFdyw
3/6qSOQR/cFmERsUYM20lnfVjfr3LW3ua04eVkclBra8DH0DLRme96Ma/zfjWh7GKnI+ZIvRYuyp
HiRfaN179wA7olzH1NWmk0DX7plLPu47sAhbqq5lZ+nblyb0ee9pIm4m8XE3ay0oxKw1DfixWnUq
fGkuc4KtDYJLM3ecAM1WQGeLKetWqnZQoQ4ZW4kvyrh6eDkVhN0xGZyVO31vUdZZjYS+GqOnzkXo
3B6CY5FrZ5JJrspUi+yrJLQBjFzGsX5eWU5H2loEKiy2p9S0ZvN7HWB+8wmZgUnNghTLc4jAIMjK
cYISX8rSCuXrtqF5zMK8THV/ik5w/oOmTT6evLFP0XvR68+KGiyMPGhbmuq855FEUkUoGoasV6du
5rbDpxWhEfhU87gTwFpfeBzvA4OV+vRJa6CYqwrhKsw8be1ysigeiK54O14QvtHBJi4Qo/e1V/vk
cUAjTpR0CWxKOZjE+XeFtZu9kbgp2Ra7iWqGHHXdq2eVbFjua5FszoLTwbxQr+LyoHLvhsZNaJG2
9r5EcoM7nKYGAqaRRZgYFy9X9UjhetANyPR38KFD8kW0NQzUpvwCLJ3ppsnietcQvJcsvdRY5YDT
CcPCaJ7Xg8rMXY/w84ya/+UndKf8yLkO8B7pxRj0orE8VgnaJo2W7RtfO0/f7+rsCDAHWxaqWiMb
J8F01drhPiB01PEGoAhKe5d3L9gAJbGHDBqvgk5x+GmvklnMWjuZyy9B4hKmLIEz2ihbM9n5GOj6
ZNavYPJPJ3ui3CniVPBva4XeKSXBivtT3oAGjQtZIZ4HTsdqFPEYu3VwUFpv+Wl3YuY9CDQ39Mq2
5j8OmZHM0BH1Dhdj3DakIB8fp5zzqJ1YOZzjVqjh94ZWUF1BTguJJMNckBbAn5zMFLgdraWKYnmB
p6OKA9bnBJDDWumEMkXlYj595nFwWU1EjUrgBN+tlFilwV86HwK1Wy5V6t1k1k8nRjhMGCkehWuj
/J4AXHrbJ3m3uJEZXyFVMQlCBTuw/7GxyQVXoIPrUX7AXCS3nZku6z+gI4/ygVOILdDfLuv8BFW2
erGhKOJqAZVLXyIm+27ML6vuaelv2E8zGRCK4n7l6RtiubGKLwWNBfkhaTJ2xPd2ew5mqJ4z/t/E
PV60Mw1V920u9XulCqAWf1CNa7XY44Vf/CJeQXI94Tj1Cm7Ni5Q0xjj82Tt0eTEkziUZcsjjON3s
I3i487xcKtNba/YWpqgpPR2PA4+plz0Py6BOC3ruCJIGPhdTm6K6tOUiQbtS/H4+PWaF9JmbobwC
RJ40r171uMWtjclO+eYQJcGAaWYwXKF99DUZBbG7d0GExX31SZctKRHPqOUvzYaNnc0I/JIswpUJ
JQYI48Ts6pp6WWsoCCSBfuhyxa75Bt8SjLwWF5FoYxvXu7zvuqxKWfaepJXelq+k//9jQqW01dCw
UFyKPBmSWJ0xrkw7+CWdaCnlsnjGn4wbhgQn8Y1Athadt0jo9aRFW3Nvdz5qK999gWT0rCUGwdnR
Lth4XK7BwbFFyYqVFOYNlohBGPyGrfjv4rD9BeKQxv7BygC7n+w7u2+G3Y7HjX0+EpbtlS0r94j6
DA8dl5abFLVP7hM2922tZnkm2GRB4+lQBJzpsQ7ANmtnDrsXHLLHlB298EVniaaAZ4E8D81B0g+v
AM0xcjAobwvV1HQSj0pSe04XACt2UUWpXYMiKLe4CoTn3xnOR7mD3+5dNdhjK8Fm96d2LArCCRqJ
QDYVwev5XcskO1yMx5MCMNC2NrG5mVmyp6/Ama5Wpd78tjE3Ysy7emqZHmmoIi7byKe40jyIoGHs
f+jTwBdUFO1aYNG/uvlKQ1KdoCv+cvkCyvvD/O0U6jwF8DRnAdHh2+OeSrKDHf3xsno0n6hT7oFu
lpLEaGGk47jUuhzHYhEbVe6wKYgf+vGtM+5D6AWrxKPvggKvJkDdFlqCBSZqZz/Sn02kJ83LTArR
fX5ORUyCoCPZk+mMMHqPg2OKN6VwZjzettFaivrhFVxWyaoyualyFjCWapLTBZLeMhd4ZZ1WhVB7
X99yuNC+uNeUMChnIE0YqyAlB1GslZO3k6IIqOlzkreNQXWzgAUuUo2deG3r9fXtXfJdbALS/orE
RgBJDxSrP+4OucKsIupVv01xPIjDHdGBYjjy4Iyt82XBnAhJLHoP8YO5sG6Bud8BgRtS16LElKga
D0tiBEQVmQSe3TTl8mfyX3v4+X5A4ZEXeIHhPXrpXQSwAqsyOBb3MlextWz6SxfsRx7Sd41OJbdK
oo9JDNspptuQPMOcQ6bq6BkFPKtEDdH6ciQD4X8jzX1Cc1003U48UmwTOlfDFAqlYfvlF2HHKS0C
Elqu+X7Xgvow/mC2L3YagbtdwzMpTwaC9ZDCiGXy7Xm9WcnELggAIgjXH7RIFZ+8SFO6M1M0Qw4+
yoNz6VPZFD+FnQBxU3ILDKoABUjas1BSn4cS72Q1I7eYMQXS0aXWzrNaZRD1ZfeMy1L2iNLcfsAh
pmle4dcmFGCC6FwYfKtU3nxO9KLmSzh1/gxJC8Vb+R7Au+dItiPWGXO7eK8Nb2P7A4+vL6YL6mRZ
Jpg88sXSqashu5AAyRXDSsHeK4aS0xNy/fjDL91jPaawrw9ZHUkynGYadJKtdArIMcrS4QbjS82I
fOdF2O1zzSPdO/Qtw24QxOERQOzq9FDRVo/789t1Aul2+8cKIRq1mmnc5BeRd7lK5Be1/Az/hTXF
nFTXVzA5vLgTFg517+Agu+Qq7GHybgJl2sUN2cN1bGwa3p5BBV4otCYwj7uaZWwEr/vRH+9M3vD/
U2OFGM3gwtTL/V4L31qrKsdxiFELMlAjfo/3Fac9Gweu6ZtDzhZ5YHGM9q+AZMHVUrkB9W9Lwmk+
6B9T8nH4wO3GQSGqVLeWfWWmgYmo9hchhCaG8wlylztqVajNd6TQf1/3dt6VwkBMfNNe4Jk4XX5k
WmX0EuF58CaEMT3zAiouwttC6sOeGYhjHM/smquyk00BfFMrO/+DSHeF1gkc5u3T4oe/BS9D9n3N
DIZ6+zFmB/Z+BSgK70NxBA9srumoQl5XVi9+IfUlyNtEVGboXWXUCBu5Q/CnsoDcTakmZuY/iPAL
A7kRl/PNDNCSwawvsAmqZKG1rXPDmbdJso2yBJdAivcelBClnUK8Zpp13Hgjn5l51PTew6MaGJ/K
SxK8teZb9uW95DF2aLawTCKCdbM+qUAFGEwdv6q7zcN0tjQIqGYAeHfKIYF3VUbTO+2lPx7/FW3f
Xs1B+UoFsclniIb+r4+IjKKYkDLJbrtOiV0N8/m47ze3yE38qOiXddeSBnBx8rlhy5l9uyUk884p
LqNWgXmKfL4QDNDnHHI4bwY0+05mvZ7NLKCAUywyxD8FDiihwnDjL0OuQdcZUyEvSKgOpv8740+C
ceK7sBhV70DYmMuBN2uLLzrlBV1MR8H2crM7ySEbe//oazLcGeunREOmqveYKn7gjUufzt2VAGdO
Mjhbmx3yzADT9rSQbUuqnYQ8hJdlfsYWVFBRGA/m7mMvRHM0gd/C/WzivSquMyr/Yt1nNIXnTdIe
LH33vIgW5GroZJo48gMjOOX/kB07/17X7mmKiRMzrbdjrTlXc/cCKW10NVKXkoT0YuArUlEd7Yf5
cJh7PypKNmExIzzbz9Z16gAxXbYTvFgHMR5bK4sDuIM1kUZW92QZBTP3NQuCoBdt+tE70mR/Srl/
i/Asf9SG1emXoBCWGMZGZ5ZE55shu/UcbAOB24Df8anu/nUtF5Nxhs10Sd2Sf6oiwCktg5WL7HGt
9yZNKJYzIOM2slPgzQ9zknU4mYWNnE+fKmdDEAOt4nNPHn6K2IyGoBLPJpH4rAjFSGmb3eto4RNv
188XKQzk01e7Pt8q1ela6GN9KdOnIAMb4RCEnWHvxYHdEgjVLa4BYBS4a/KzOGbK/onVe1FfMnIZ
A53+dCMWalnE4H5TCPzsedyLoDWfw9g7P4TBR/PBD/ZrmkbNNnW1BXzLO4fxNqDZDHB+OHMjD5z3
4Va3zhcKGWWhtsXPJoyuS2WOFS8qXseTXPsBYffR6ncsed8K8aIEPkoBdvJhH1NKMyeH5dVif1+/
Vx/AtpuxR81jU6163DQZ0TfZCqXOgYrh0MULMP0pgQH4NqVQXMlyKusgcaKgetF8eraWWV2HSXTT
kXVFg9JPNH4cjGJibTzCjXMpJMWybV+Z/RWhifMCwbA6AEfo0W1IsDKMcUl5JXb3TZSpT9t6VqU2
hxezdeo5JD8kQ3J7tbJfXr+0PzQPWOCV5BniUGh3RSJ2pBPIrxmqRUnuupHqtlpIAsxdEM811U1O
MWpB/Wihq5/dXRmi4GlIPYKZ9/evk/SyOlFyikb5CC2A3gL2yXgSScM+wf9sXlwOFUWhedXYvGLp
Lbkxgj7MkLPrj1LMoZ3I7E8dc90aIUjzxVsXO+CvkiypornJkudwS/xueibIwF0TLwJAbxbXvUhO
5Cyl2gHULhZHLMaR6xP0SBZwCn+0e41OiKv7AJaX+ICydAI3Z+S9s6HLpz/tF9CkSJPCunVp7Txu
AP2Lw9yt/2iq6PZF0x85sKtVH05/eq2WDIMXnYPuRf7BgZWXHDbdoz2tZWGLSQYArCFhbowu4YdO
FV8t3H/fz217RtwVlNGWDc9wonJCXewWEKOG2RPaJ5Cj5KGUz66mwhLqmdPL/xgKD/CBUNjsXyrC
Lk/RjuJWuNdW2Pipegfp4eozhQ0AbCpOZlJu0wY03fTjttFYSHgfQp9SkN4Y53j3mAly5qdDlGPT
DHKHw3HaK2t/e9ksaH74Un5w1gLX9vFEAz0guGaKv5/MtM5oHssUj3W2Wg8cDjJ1cevxUeOjPTqG
OfSi5K9DuNDVcMJH24JNqDxrU/LH1nbsH3AIeelds6sEYvvS+q0HptvadyLFcTxJBfBZKzyucy0A
TL8QX7BcCaMo1rfnCQFersY+wVyIwtzeTY8OInlIVSphg9pf4fHNI6FRawWa2IP8k/NeB7Truvjc
PGAX5fhPEFzcJt9vdIYSqqSqAtLpf9sT4GgeoQeastcwiefSuAW90tdgRpzgjuyBx+CxrSgtXiqw
MyWCi6THtdwc2oNUcV++aI4BN4omyg6NUD5I+enGO3mQ3zPARppEzp4q5DU802/08B8gFPHNlAfL
3de0mH5LBJFYggfftoSkZnWgcbERPd63R3ewP/PaHG50Q//QS2iNOIsbL1iHtK6wNnrdLBEo6N1r
UkUMn/4dHynyJuUUdODRtrwfawayN5z/ZnJi3RL1+ZPJfFqmoGiuFixGrVUEuVXEGL2NdbRooJpC
vTUgI463+ABh8uXLQlZDhtOd2yvvaQ480KvENW9HvFYjBkRw2T/rL4hFbEpjGR8guy/OY/HihmCx
09NlJCftjc76HplmWDEsEmUjpIs59HnKnBGYYZLXzqW1hWzJwlCcZaUvS3Km1uX2o+oyzAHUAoNG
XgOCdFxlJdyAcfgOFMiEVX7J13K6W4vz9DB5bZIh+NpwrUyRtK/qiT/xkjvyv8IcGgAgMgZ+Tsdw
nrAdk+j0r7SlA1v6cTraaeNwZ0uHTUk2UluG7MzvJUYHw6lI90WmHWrPxB4BnuWZaDBiHLSgAXVF
BTNMN6+5S2M9hqbeJgdg7pHiS5ZvoGLjdccvN7pjvSvOyeh1hqSyMXqxIo7MQFU7gdYKs1npe7c3
S4lwYVkXD4eCd54MLrDrR5/Q1RqgOcq3fcx1FcYvz8gaF0fdABEaaA8jq5XnZAyXDp9LmeHSMa7c
LhXvE+IDe5K/CCoLVrn8Kt27uwAFUzbP3FkceLCWVkUd983Cdivkce8nbDOYPe3/9/WaJEvD15Pn
o8vWtm5BbCE6eILK7GV7jz47b8E8Iz5CYo3Iuc3bIuuz3E2IVFRTLfhzmH/Mib6WgcIAitD9nVGu
U560pgH6thAv4tXqJ/mNMLZwP4rPzdkSTR6gJZNxKE7RROxTPhofqlDQGuCHodU87+Ojs3Cdf66h
Meo7BNtLVosk1XMMk04t4ptREdTWZs9Z0S/w37db2pXe07Yjfeuq2wQdFDRlaIBmUDf5MADHVzdO
SoRBpEkGxEIOUV5i4n8XMlDUJcqAkTJTGxJgT47gH+CqDfrpnavaAa3qR0JjI1IAMioEHg9fBlqx
7dunZSG1oZ/hDwVURKOXD26KpyelKLSiHzPWNdP+iNc7zRAOOahOVXMO+eteyh40QrKmZUM/dp7j
v047nTqFji2b/Yc2sLoHxagn8x8K7r8z0gM1pQVdp+cBxgxXpMwsh7LjnQpglpiHp6xMKRr6Tg1X
vw6/nrl3bnMVJqMTzoiZC8iYj4ESjVatvO4DRaEceUemqE302HUZbZj9tLZlhWqpompoaBv2YE0+
GKb/dBFce7oi1ACzSXh0UNzr293X6+rOJVJU2TQYYbRHOklOQ+ec1KhVO0TTpageFVO3y+ymNmXr
y3Err/CtBbEga1SJhjQ92JDp3hUoDEh6dwtmw+GMkQQxu4SymF0OmoERMX+UhlLZKt3tUOngxoec
sVJpBNAuPDjALmRkeu0Uo5M8HEFLN3TOjP+vUbQ1RqBDuK+SukkGg2yJQW1q/xF6L4nTeRsksaNn
pbLKDTasbchzWtc6QA2KyYu7ez4rx53CRkCFHt18NQTm0QPE8Y2j8MJm8y3rbaPa60TKD3kxwNVb
gf4KRG71lQnU9YT16c4MB4UfM1L3p3/t+vM+21Lk3dZqpzbVOmFSvUli8x4g9yKGiRmjoJ5jl8ni
PGFimjzw3aKx9qEntDEW7AT/ejPN7amP0AN3IrwWINPK+2wvWgLjzpf8HB/SCscjcf0cY8qhHwk6
/Lcb+34vK0tEAashZPAwGe3uzVa1C9+CV1d2ZmdrCOijhEIGBM8KatmBWMTpx5/o8mLHtsvQJ49S
8FFEJkfKV5/KHGQQkiPpRby/LcauKfEoma/Tli4FmpsnLAOfUOdr/7IJ27ZYlPnrmNV29E5xo6TZ
sOYGxnzAAHrfEIjj26RBtj4sNLlG0HZ60iUIkZUHYQ387ppLzss0JpjHZu7qWBouSAiLkopoU26n
4Qy4O5hhq7g8xnsCQ39HiiyRiMDvX0u1SuAAFp1UiinI3SsidfLZrlYuUgP4ism7g4zhIMrAU5lK
+NB0j0kSYIAHrOn7Qm9SVJGGC87LJEgim3N0FiWXOkkzRWPpSKss48vlc2hSsPEp0K5Y8VWxHSzi
b+IODRw0+/z1L6Z+GS3lKvnX88zqKWYxg/OhsN4nTg6MjGIx825ZNMMeqHAGmFQQFUC5r6UMVrXQ
5TT0MBC2ZHDGVw0dpy7E7eMn0IAnSj+gA0qdOrJq8Wievq5K8lkUTeaCEqoln5DQ0JQVRvvhu4Pr
WRz7rE8gtAoVv79HRFVbPhDf/o4NQz6A6giuduWrU6Tqj0WtIFPvzTOT2/aB0Skt8Y6J3zOlLjNO
CIecN2/SAI+v336eB+IeL5kbNK80A1yRi0SIJ798/6WiOFPtdCGO80n3KKpmEx6prc6IopEXXYI6
dLe6motTFnfUkOFy66NMDScXSLbE3NKMDLVbGItvtkH9O1NmLkyQHJM8Uw5gBM6vE7M4bN/7uIfp
WHVlBhhEYfV73LHGYZuiCp7pYXLNXJRTZdaAwTdCDtDJOILFdBGE2OcIksq0u4ZKb8E54QEI8hO5
kjlXl7KT7vJNyaYCJ4k0BGzJ8pnsgXBRWo4IcAPqjXyXcVj7YWmbdK1uGaBO51ygEQaACZyKj+J5
UWZX2dbIwceOp5zd7EsDbM4dXcMmwXZ9ao5tjXmY/VGId+plQEy1eg/++Ic91G1qsozMA4kEq4lH
hVk7v30F6wQEE8FgWOvEzvSQlvDRLCinJzW6J1+L1KzT3dJuz1TBd1aT2Y+MVH0qJo9j0RInM1+8
CUD0tb6Otsci0tMWJFPhUacKCeU2GO9x39D7zuwrj9lo6kJyPvRkTA9z0ruHx8pBeRWlLavqXOwp
povYWeLtuDEvQajDAKu+8K0BJpKGTQxKjoHPHBQ4yBICiOqKTlqb4AUlcZEzOW0U/cjv91IPvsdh
JtVQpY5YMrwxS9D1TgRd+zUqLt5b5TJ9HE5JdPrNSvGYWsf2vKFLs8rnF6Zw0nJE0JzXXgQ2x5jl
qYyaQhTF3N8kPJO/Cc5EOlzb/U2OAnaOW3uKq977FQIzLoS/5cowHadSiGeDQloFwdjMghkkKlbS
oCLZJK+smCXd6/lnK9w9/VQiCYKMp3JKGB2OOWuIJ0yTqpaKjPNi+tyzb3fGuScaQy1eH84H5iPC
gXHugkK0GTMBPuphPBDekIFBH72W7Q3S8AVzwFNyX/jFF45ftokGx4Ox7o0y7k/7S+1p5JBrUioF
wrxrq7v467laWf+o3InIRdXZ/msJm/ViRVUkXsRL/qUU/V6bLPBx4oEPUnntZYUtkjf9W8in4aZ9
ztG9q8oGuj+L8W6jVm3pusDQUKACwLK22rWmlmqsV0mxfOtZsuW6siLe7lgyYZG57Q4vUTU4FyR5
cGYqBsi3d2U/eqNLmEwV1PLpUyX/1duUkH4SjUOQ2/F3RgO874OpARV5jGYAHalVnEXXl/Jwj/F7
t8fUEHI9vAF7PjbMQZj602FvxE+5mpUKHxhsx8jr6llZbRWkQzInlxikIhv75qffrX5v8hEj1/SO
OzORtC+GLENWvu4M+cUFf2oyQt552uyLdKNjK1YsnsR003Nes91dcKs3XzMrCewjtRR4MuE8B4A5
HJtLSHt8tAoZdMTd5rm6IPSoQRDuPSLlrSOI1Nrf3qwkZ+y/oy9TxpvKgcKC5EsOiBveT38oQRr2
fEMB5NEAv39YUOd/MrwBJLzqcyzHOvZmG1xTDl9DD/gfR+WsjvkrakEdMhVLnJfLY2wZVdLlx/Tm
WaimlBrA2ufXmCMIcsZS7H+4JMALPsoPJPBW0xJ7ifkKanedX3P60VgqJJzQv13BoPY982c3nDPW
G8d4xLhTQuD11qYdZsPuNntYPEU7BzRi0Smkq8ft5Et9BYIa39PrEbnSzPbm1hMcFUpssPIcGOSu
a/Zf/kwWnpoWZVjcB/cN8WNVedze1OEJ7tXR9isiLDZTIXFIsYL+BeixKzKczNJXIylL0QC1I4vC
+KqzdnkySbpVxCYlEPvbhFGF80aSxLBjRsZt5aRZgRE1JvJxvRyj3F/fmdhqsuVxXjU+1ZxUar3t
MOwoY5tLYEMbAc+DpqFcXKzSvN/wKdM5xMJhJD1X4SGwe+Y59dh6D6dUkzoVl4b8RbNQfoPwr81h
xoUXm4pWI7N6YZP0OLD0eUoqzD1BSrUSr5qhYYm0KcdVsGLHqV8CG6QvHSK1rTU5i6gWPGJaVqi4
+47/xl6WK40AuqqOMmhPZU1Nu4i8yovQC2Fc4p0D7pPR2ftMKdRuiAqtV+4aAC93duGgsnY+R+7Z
9TSnG/Ne1GSNqKv+WM0G1xynuIWKUVwxnWp9ZJ5rRUmwAiMI+N0Wmua3w+XO9vXgEmdcohKeV3uq
8iiaFUhudTIF1YGJVq6hHGJJpftWPQDLbs4p20fEdeU8IRL8uGJmAc6pezEG8MHa/ZEfrH+5vnHk
r7NPMHF5pT7Qw16SfT3ehLlZxBBzhG6thTUwrnm3cC+e7FyAvvLhMWrQRP6gLeHyE2t8CYg94973
AFHO5VZBOljFRdbWGqPEn8mBbMGz5ojkq5ak29v63fFJbU7jfkjnbHzgaVPDVSlY6Q5a5WQ2/7cg
j7Fz87sv0XOHtZZGale7x7DHbbakqZ8fiGSD7Ve+GmDeEW4bB8SX3DVnR0zYJKHEikq29H8cywX4
4FEBNX7P/xKX8Nioeq+fcbWHGksqb/BSC7dLlUfGxz+4f9g5x6lW+i2HS26oJCg+4Gt8budj3E1N
wwz6ZcuGPuJxQvh5q8iOS8reizu2t582MU/tZvSLy20dWn2b9OXy3J9Blt/kS3A0Dshx/cMkURtM
rHSBpYqWVooicx1Q0j8Rk8d/ZsME5ROk3sBbWOjG653p2+5IigYdv21suLI/Y6+asqvwhrIZq2eP
JLVjO1AM1e5Gd/8BCGz/MGF9wUl9dCNTjALUMGyld4zOrG91GNypGxbYTV7eExvD2cBiB09Q5ESp
0daWgR5xEw4+kqrp39vz1wMv+lsajQWJUF6CwiosrJfvTB2ZJ2ZYiVUy3lokpdezKFy8+dEAGCjg
VN04HLZy2Knqvh5aSI2MtP3mYre8dJbVmYuavg+GbsXEczqZ86DhRIAAvgEBwiJV3gNss/pbR2oU
OqPvYbiXzm3R8CYNGoMlGxfpTnO8r2zZH7+/9UjmYOddNpCLBoKjG3Q8X/Y9eH1fySu5M5ZVzRdO
pVzKasCAScCZQZtNqNflXlfL/B2mzJA1LcS3vhyFD9ztMUAi4SLswKM1gN7ascaTdCHvrjGRQkQ/
YfRQFWNvkpW1MUo+lbWtVtjkDoF70NOu41/HlQo2eh460A5jZhBfCT2NoSk8EkZup1m74AXA5p6f
rNBknrd3ilrkpD+cwc+JgjiKg9AFniIO9/G19tORsWR4k9vBpOtHEGhoKxwJc5b2JPTL2M+PiosZ
EU37EC17cMSCYoezYyk6T+acjKwq/9gk5+bFIQ6C5ntvkzgsPxvhEyPsnETHmeamtTVLndoKOYsd
KSUhYcZiAm351MlQ416Y/Mofi5QB2xCB+0qah7kly+gvyNNSNXCDDXYRq/lO4f9WYM5Bc3+XWgNd
5Bg3sYkAj9luEuQ/d6dcmSqVchdFTqME8CtJsuWlvNu225ZfRU5TxTHlCfINn2kzPHJPIFq9XWkR
c05e1NKvACD4ND3+glnP9yOmQdOpR190ZZptVCwjjE91mBNPWqnm683zlBWLhc33hVgv7CL21HJn
/yBnGfTjziiUGgyWlO3n9pVkBgVVZRJSQrVIwgixvIQ7k9InbuS1dgctG1xlMn3ixEArXAusstiU
U7X3y1MA3zEkpKXduUjblYxSpdI7LpiFvJNQ2DQ85SmgLQHFhycoHDdpWyj0MY4OQVGXUcTU77DQ
uT9FUANAFV5dACv/IVUOD80ilNl+SxLsBgIL6RVAsL03I13gnpWcCMj6XBSUKCZKdEtQIkhLpayt
fGD7JQyIbaMJ9xxfD7tlFs+97DW0/ABRIi6K0MTQW/w7eey6nsR/AFWrQ8lU4p58hvz17rbQSuQf
FAgGECi4qw9/UdNr73rOHtvfWhK4cMR9jyChs9dto6YgFaUUpxWMIVgq1W+QtNoHTxq/cQUT/tYu
nFNS+uZks2LZe2khik4OaJnsf7jivhIQrbDrQaMiOKyH69z9Vu20UIFDU2zx54IGTP5S6OiIilVE
gAUVVAmgIYpFXWDjuURvmXuWB6Zfx3zKadXi4xnaNuATNWrJLCcViXmDPl3tPnoHxKSvatzf8ANg
oYdQ/0LRA93egKV/79H1XXAa062bX+Xd0wRGnljDSbJf6XUp/EqHCvSxkha4AthJOuqDk03zfuc1
n5KCvRTnFKWJ+YdF2szrq0umBKfVQXts3H+upPltG1klpMsxTf0seP7VwVAthTKezE6XvWHVgm/q
oGRBy8xnNa2gBt8e6qJtMHeC1xUQrabOV9a1dqWZaPV9lD7dLuOousp/I9JMdYeDKA/wjC4wpnE6
hMhi88y57K149+fLmcr5OyBLcrbso6iATiFeb1xG8OyrQE0+e5ItaG/u59BwSkvse5fF7Rl01lR5
XqZYymK58ri+Am2jMKXI0nlozF7YUj0FK5h5QECjdznLeOQAbvc6vT1Y2lsgPv6jnpTJaKlUUHZz
ghSXWqXeaUH5moXemCp2G7Sc40y8TS8Tny3evtESs1vM8ATKZStq/YkM0HNzevHiZWj43AEBHzl7
lt4ctNt0uBUrUQTRSByRhDKHqRKMPr28MX5g5dWBt8fXjdKBKYq/dXrd1QQE+G/6SQYN7TWUEZbq
0ei2JyPIKQziINxS7IZpzR1jDND/H/gw1O7bPtRjEuToaY4HXE9uX7h13vRX0Ahg4GUUCzllf65g
ES13PqRLz6be2A2rpIhaGuklEV/6saXsoXGbg0Ll9G0XEjGIQLa1f1Omq/DFnaAQIp42t/Bp5Jvd
4A7OWsTTpywbY6e8wZcfT438AbyARvkT9szTrKDY3YMcmWjpjsVdZUZ9FDV2kHzrOtLyEYcC0/rZ
pH1fLJ++IxldxzpyiSRIKIC0oHeDlO+oNPM4gsH4B0UH+vJpn4ZiGiTZVRcbVkb+e1cPXNR+pbcI
0kWdIiIUWb+EOg6NmzY4Or5YtzlRe7krQBGglfmTNtMy6aUFDTe4bF2bUieB4Ay0M++dGi0989MB
UsuCFcZUWv1m1K/BxD19GUCatJ/d3XsvosX5ahVNcw41TXkto2PPdCobY20YO8SIhyILQt+68CQQ
2nYD+9oT8FCrtthwWjDlzfRAgpbZv/OzRxk9zJwSu17NZtmxh0j4SJS6OaLN+LwyxrD9SDBSczWg
WkW9QkgjSAUX80JYR6Ptoo8Pk1EIx17uu3SeOhK6LFVSDuDLXl9tQxawbv1Dfcq4Xt0sBQBZUCAX
k6/tVikZcYRwtf33s85wsjXaVKzApgYoIKgrV+gP9aaUiTD5QN75okkDIPDzjK3jlCNNgXUWirBi
AqfkAVWnjweoBfj8lZDAv4OhmR6LDZLN1m398BI8BeXiCrCIKDLV9Pa1RC/LP6soB35IpbydUhDK
sX5aGOszEbHqsXKd2b7Iv2QwX7U4tMDlBc1Ull036opI9LujyByffeEUQrhEzmMFGBlcpyyi37S3
9HcYc5NePXi/9BTdwOLRJNgb88nbpHH2L+Fmm46p6lVeVEtb5TfXeUU+gLGS0hHLIPkcx58t8VHW
aUd6wqjXC6FcH7IP+k7tcHPiOjE51VH0kn5OPfkc9JpC7vqtcevtud5YgJduSA5R2KeOz7H2llgD
3xCJgpOrsDuhe/FT/SHxhevhySRU866n1Azv+3Vvi70zRn8e83lHWnko4rBgkguJOOiFsW/Gs4fN
z2zGAP3M7+On9lyVtnj601MWfxvNJqXm+lPEYrocw4u2GMlrCw+iZlBk+ZXtBAd+b3HjzQ4FF9HH
eTYwka7nyQILqsmFE/6tWNe194YrXSG2WK/Gr6Xlen4dEAhhcbC8A+xyy3dasBdeAp4W7XU3p8/Y
uRpN9B1NyVEL2uqp99pKccAdAo+pAwtq3DSHjTOQrshQ7wd/arGrXB8xFSq81O640d4eIF1Vw1p3
0JwSgZu+JmW2R090r5JTRlos8/+CQnEggOhthlrUhG7wuJyKI5i4JjQGN/HZ3G5VGggtiA3th8W6
WcHzgE6fdvUiJH2mjdmLpEhySw0NaigQNFQY+GgNTiViKQVBBnKZmMEK9sfdbl1zq346I2xnLId4
Q9GyySEik4sS7EzM2e8zvB690P1AsGyqnYC4DaZ/7zhtTGFwzXzKkyoEkoEH8LMcaOnzHeqwTp5J
ECJagIB5b1+2olqAYoq0qHN6uEpfCIKcHSmJdCaLNFakkt1mKGFVyc0VNpm2My/cOrqBsEQHLbLR
YFM4Kr6O4Z90oOxwBkyh6JvAUnXerFZrty2dT+f7GbKMqF4IKj/GAGAf0Mx2AGRFzgZbH8bRMaix
VI6zg1qqy8Hl1Axg0saU50oyYg==
`protect end_protected

